// File vhdl/fpround_fpround.vhd translated with vhd2vl v3.0 VHDL to Verilog RTL translator
// vhd2vl settings:
//  * Verilog Module Declaration Style: 2001

// vhd2vl is Free (libre) Software:
//   Copyright (C) 2001 Vincenzo Liguori - Ocean Logic Pty Ltd
//     http://www.ocean-logic.com
//   Modifications Copyright (C) 2006 Mark Gonzales - PMC Sierra Inc
//   Modifications (C) 2010 Shankar Giri
//   Modifications Copyright (C) 2002-2017 Larry Doolittle
//     http://doolittle.icarus.com/~larry/vhd2vl/
//   Modifications (C) 2017 Rodrigo A. Melo
//
//   vhd2vl comes with ABSOLUTELY NO WARRANTY.  Always check the resulting
//   Verilog for correctness, ideally with a formal verification tool.
//
//   You are welcome to redistribute vhd2vl under certain conditions.
//   See the license (GPLv2) file included with the source for details.

// The result of translation follows.  Its copyright status should be
// considered unchanged from the original VHDL.

//
// VHDL Architecture HAVOC.FPround.FPround
//
// Created:
//          by - Guillermo
//          at - ITESM, 11:08:16 07/16/03
//
// Generated by Mentor Graphics' HDL Designer(TM) 2002.1b (Build 7)
//
// hds interface_start
// no timescale needed

module FPround(
input wire [SIG_width - 1:0] SIG_in,
input wire [7:0] EXP_in,
output reg [SIG_width - 1:0] SIG_out,
output wire [7:0] EXP_out
);

parameter [31:0] SIG_width=28;


// Declarations

// hds interface_end

  assign EXP_out = EXP_in;
  always @(SIG_in) begin
    //   IF ((SIG_in(2)='0') OR ((SIG_in(3)='0') AND (SIG_in(1)='0') AND (SIG_in(0)='0'))) THEN
    //   IF ((SIG_in(2)='0') OR ((SIG_in(3)='0') AND (SIG_in(2)='1') AND (SIG_in(1)='0') AND (SIG_in(0)='0'))) THEN
    if((SIG_in[2] == 1'b0)) begin
      SIG_out <= SIG_in;
    end
    else begin
      SIG_out <= {SIG_in[SIG_width - 1:3] + 1,3'b000};
    end
  end


endmodule
