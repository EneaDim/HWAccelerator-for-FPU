LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

entity tb_MBE is
end tb_MBE;



ARCHITECTURE bdf_type OF tb_MBE IS 



COMPONENT MBE is
    Port ( A, B: in std_logic_vector(31 downto 0);
			P: out std_logic_vector(63 downto 0));
end component;

signal Atb, Btb  :  STD_LOGIC_VECTOR(31 downto 0) ;

signal Pout_tb  :  STD_LOGIC_VECTOR(63 downto 0) ;

begin

uut: MBE PORT MAP (A=>Atb, B=>Btb, P=>Pout_tb);

process
begin

wait for 400 ns;
Atb<="00000000000000000000000000000000";
Btb<="00111110100111100011011101111010";

wait for 400 ns;
Atb<="00100101101000000000000000000010";
Btb<="00111111010011110001101110111101";

wait for 400 ns;
Atb<="00100101010000000000000000000011";
Btb<="00111111100000000000000000000000";

wait for 400 ns;
Atb<="10100101111000000000000000000010";
Btb<="00111111010011110001101110111101";

wait for 400 ns;
Atb<="10100110100100000000000000000000";
Btb<="00111110100111100011011101111010";


wait for 400 ns;
Atb<="11111111111111111111111111111111";
Btb<="01101011010110110110101101011011";

wait for 400 ns;
Atb<="11111111111111111111111111111111";
Btb<="01101011010110110110101101011111";

wait for 400 ns;
Atb<="01111111111111111111111111111111";
Btb<="01001011010110110110101101011011";

wait for 400 ns;

Atb<="01000000000000000000000000001000";
Btb<="10010100000000000000000000011010";

wait for 400 ns;

Atb<="00000100100001000010000100000000";
Btb<="10110000100101000110001001101110";

wait for 400 ns;

Atb<="00000100100001000010000100000000";
Btb<="10110000100101000110001001111110";

wait for 400 ns;

Atb<="00000100100001000010000100000000";
Btb<="10110000100101000110001011111110";

end process;

END bdf_type;
