library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use ieee.numeric_std.all;

entity DaddaTree is
generic(N: integer:= 64);
    Port ( IN1 : in  STD_LOGIC_VECTOR (N-1 downto 0) ;
           IN2 : in  STD_LOGIC_VECTOR (N-1 downto 0) ;
           IN3 : in  STD_LOGIC_VECTOR (N-1 downto 0) ;
           IN4 : in  STD_LOGIC_VECTOR (N-1 downto 0) ;
           IN5 : in  STD_LOGIC_VECTOR (N-1 downto 0) ;
           IN6 : in  STD_LOGIC_VECTOR (N-1 downto 0) ;
           IN7 : in  STD_LOGIC_VECTOR (N-1 downto 0) ;
           IN8 : in  STD_LOGIC_VECTOR (N-1 downto 0) ;
           IN9 : in  STD_LOGIC_VECTOR (N-1 downto 0) ;
           IN10 : in  STD_LOGIC_VECTOR (N-1 downto 0) ;
           IN11 : in  STD_LOGIC_VECTOR (N-1 downto 0) ;
           IN12 : in  STD_LOGIC_VECTOR (N-1 downto 0) ;
           IN13 : in  STD_LOGIC_VECTOR (N-1 downto 0) ;
           IN14 : in  STD_LOGIC_VECTOR (N-1 downto 0) ;
           IN15 : in  STD_LOGIC_VECTOR (N-1 downto 0) ;
           IN16 : in  STD_LOGIC_VECTOR (N-1 downto 0) ;
           IN17 : in  STD_LOGIC_VECTOR (N-1 downto 0) ;
           P1  : out STD_LOGIC_VECTOR (N-1 downto 0);
	   P2  : out STD_LOGIC_VECTOR (N-1 downto 0));
end DaddaTree;

architecture Behavioral of DaddaTree is
  
  component FA is
    PORT(A : in STD_LOGIC;
         B : in STD_LOGIC;
         Cin : in STD_LOGIC;
         S : out STD_LOGIC;
         Cout : out STD_LOGIC);
    end component;

    component HA is
    PORT(A : in STD_LOGIC;
         B : in STD_LOGIC;
         S : out STD_LOGIC;
         Cout : out STD_LOGIC);
    end component;
  
signal outpp0L17,outpp1L17,outpp2L17,outpp3L17,outpp4L17,outpp5L17,outpp6L17,outpp7L17,outpp8L17,outpp9L17,outpp10L17,outpp11L17,outpp12L17,outpp13L17,outpp14L17,outpp15L17,outpp16L17: std_logic_vector(63 downto 0);
signal outpp0L13,outpp1L13,outpp2L13,outpp3L13,outpp4L13,outpp5L13,outpp6L13,outpp7L13,outpp8L13,outpp9L13,outpp10L13,outpp11L13,outpp12L13: std_logic_vector(63 downto 0);
signal outpp0L9,outpp1L9,outpp2L9,outpp3L9,outpp4L9,outpp5L9,outpp6L9,outpp7L9,outpp8L9: std_logic_vector(63 downto 0);
signal outpp0L6,outpp1L6,outpp2L6,outpp3L6,outpp4L6,outpp5L6: std_logic_vector(63 downto 0);
signal outpp0L4,outpp1L4,outpp2L4,outpp3L4: std_logic_vector(63 downto 0);
signal outpp0L3,outpp1L3,outpp2L3: std_logic_vector(63 downto 0);
signal outpp0L2: std_logic_vector(64 downto 0);
signal outpp1L2: std_logic_vector(63 downto 0);
begin
outpp0L17<=IN1;
outpp1L17<=IN2;
outpp2L17<=IN3;
outpp3L17<=IN4;
outpp4L17<=IN5;
outpp5L17<=IN6;
outpp6L17<=IN7;
outpp7L17<=IN8;
outpp8L17<=IN9;
outpp9L17<=IN10;
outpp10L17<=IN11;
outpp11L17<=IN12;
outpp12L17<=IN13;
outpp13L17<=IN14;
outpp14L17<=IN15;
outpp15L17<=IN16;
outpp16L17<=IN17;
outpp0L13(0)<=outpp0L17(0);
outpp1L13(0)<=outpp1L17(0);
outpp2L13(0)<=outpp2L17(0);
outpp3L13(0)<=outpp3L17(0);
outpp4L13(0)<=outpp4L17(0);
outpp5L13(0)<=outpp5L17(0);
outpp6L13(0)<=outpp6L17(0);
outpp7L13(0)<=outpp7L17(0);
outpp8L13(0)<=outpp8L17(0);
outpp9L13(0)<=outpp9L17(0);
outpp10L13(0)<=outpp10L17(0);
outpp11L13(0)<=outpp11L17(0);
outpp12L13(0)<=outpp12L17(0);
outpp0L13(1)<=outpp0L17(1);
outpp1L13(1)<=outpp1L17(1);
outpp2L13(1)<=outpp2L17(1);
outpp3L13(1)<=outpp3L17(1);
outpp4L13(1)<=outpp4L17(1);
outpp5L13(1)<=outpp5L17(1);
outpp6L13(1)<=outpp6L17(1);
outpp7L13(1)<=outpp7L17(1);
outpp8L13(1)<=outpp8L17(1);
outpp9L13(1)<=outpp9L17(1);
outpp10L13(1)<=outpp10L17(1);
outpp11L13(1)<=outpp11L17(1);
outpp12L13(1)<=outpp12L17(1);
outpp0L13(2)<=outpp0L17(2);
outpp1L13(2)<=outpp1L17(2);
outpp2L13(2)<=outpp2L17(2);
outpp3L13(2)<=outpp3L17(2);
outpp4L13(2)<=outpp4L17(2);
outpp5L13(2)<=outpp5L17(2);
outpp6L13(2)<=outpp6L17(2);
outpp7L13(2)<=outpp7L17(2);
outpp8L13(2)<=outpp8L17(2);
outpp9L13(2)<=outpp9L17(2);
outpp10L13(2)<=outpp10L17(2);
outpp11L13(2)<=outpp11L17(2);
outpp12L13(2)<=outpp12L17(2);
outpp0L13(3)<=outpp0L17(3);
outpp1L13(3)<=outpp1L17(3);
outpp2L13(3)<=outpp2L17(3);
outpp3L13(3)<=outpp3L17(3);
outpp4L13(3)<=outpp4L17(3);
outpp5L13(3)<=outpp5L17(3);
outpp6L13(3)<=outpp6L17(3);
outpp7L13(3)<=outpp7L17(3);
outpp8L13(3)<=outpp8L17(3);
outpp9L13(3)<=outpp9L17(3);
outpp10L13(3)<=outpp10L17(3);
outpp11L13(3)<=outpp11L17(3);
outpp12L13(3)<=outpp12L17(3);
outpp0L13(4)<=outpp0L17(4);
outpp1L13(4)<=outpp1L17(4);
outpp2L13(4)<=outpp2L17(4);
outpp3L13(4)<=outpp3L17(4);
outpp4L13(4)<=outpp4L17(4);
outpp5L13(4)<=outpp5L17(4);
outpp6L13(4)<=outpp6L17(4);
outpp7L13(4)<=outpp7L17(4);
outpp8L13(4)<=outpp8L17(4);
outpp9L13(4)<=outpp9L17(4);
outpp10L13(4)<=outpp10L17(4);
outpp11L13(4)<=outpp11L17(4);
outpp12L13(4)<=outpp12L17(4);
outpp0L13(5)<=outpp0L17(5);
outpp1L13(5)<=outpp1L17(5);
outpp2L13(5)<=outpp2L17(5);
outpp3L13(5)<=outpp3L17(5);
outpp4L13(5)<=outpp4L17(5);
outpp5L13(5)<=outpp5L17(5);
outpp6L13(5)<=outpp6L17(5);
outpp7L13(5)<=outpp7L17(5);
outpp8L13(5)<=outpp8L17(5);
outpp9L13(5)<=outpp9L17(5);
outpp10L13(5)<=outpp10L17(5);
outpp11L13(5)<=outpp11L17(5);
outpp12L13(5)<=outpp12L17(5);
outpp0L13(6)<=outpp0L17(6);
outpp1L13(6)<=outpp1L17(6);
outpp2L13(6)<=outpp2L17(6);
outpp3L13(6)<=outpp3L17(6);
outpp4L13(6)<=outpp4L17(6);
outpp5L13(6)<=outpp5L17(6);
outpp6L13(6)<=outpp6L17(6);
outpp7L13(6)<=outpp7L17(6);
outpp8L13(6)<=outpp8L17(6);
outpp9L13(6)<=outpp9L17(6);
outpp10L13(6)<=outpp10L17(6);
outpp11L13(6)<=outpp11L17(6);
outpp12L13(6)<=outpp12L17(6);
outpp0L13(7)<=outpp0L17(7);
outpp1L13(7)<=outpp1L17(7);
outpp2L13(7)<=outpp2L17(7);
outpp3L13(7)<=outpp3L17(7);
outpp4L13(7)<=outpp4L17(7);
outpp5L13(7)<=outpp5L17(7);
outpp6L13(7)<=outpp6L17(7);
outpp7L13(7)<=outpp7L17(7);
outpp8L13(7)<=outpp8L17(7);
outpp9L13(7)<=outpp9L17(7);
outpp10L13(7)<=outpp10L17(7);
outpp11L13(7)<=outpp11L17(7);
outpp12L13(7)<=outpp12L17(7);
outpp0L13(8)<=outpp0L17(8);
outpp1L13(8)<=outpp1L17(8);
outpp2L13(8)<=outpp2L17(8);
outpp3L13(8)<=outpp3L17(8);
outpp4L13(8)<=outpp4L17(8);
outpp5L13(8)<=outpp5L17(8);
outpp6L13(8)<=outpp6L17(8);
outpp7L13(8)<=outpp7L17(8);
outpp8L13(8)<=outpp8L17(8);
outpp9L13(8)<=outpp9L17(8);
outpp10L13(8)<=outpp10L17(8);
outpp11L13(8)<=outpp11L17(8);
outpp12L13(8)<=outpp12L17(8);
outpp0L13(9)<=outpp0L17(9);
outpp1L13(9)<=outpp1L17(9);
outpp2L13(9)<=outpp2L17(9);
outpp3L13(9)<=outpp3L17(9);
outpp4L13(9)<=outpp4L17(9);
outpp5L13(9)<=outpp5L17(9);
outpp6L13(9)<=outpp6L17(9);
outpp7L13(9)<=outpp7L17(9);
outpp8L13(9)<=outpp8L17(9);
outpp9L13(9)<=outpp9L17(9);
outpp10L13(9)<=outpp10L17(9);
outpp11L13(9)<=outpp11L17(9);
outpp12L13(9)<=outpp12L17(9);
outpp0L13(10)<=outpp0L17(10);
outpp1L13(10)<=outpp1L17(10);
outpp2L13(10)<=outpp2L17(10);
outpp3L13(10)<=outpp3L17(10);
outpp4L13(10)<=outpp4L17(10);
outpp5L13(10)<=outpp5L17(10);
outpp6L13(10)<=outpp6L17(10);
outpp7L13(10)<=outpp7L17(10);
outpp8L13(10)<=outpp8L17(10);
outpp9L13(10)<=outpp9L17(10);
outpp10L13(10)<=outpp10L17(10);
outpp11L13(10)<=outpp11L17(10);
outpp12L13(10)<=outpp12L17(10);
outpp0L13(11)<=outpp0L17(11);
outpp1L13(11)<=outpp1L17(11);
outpp2L13(11)<=outpp2L17(11);
outpp3L13(11)<=outpp3L17(11);
outpp4L13(11)<=outpp4L17(11);
outpp5L13(11)<=outpp5L17(11);
outpp6L13(11)<=outpp6L17(11);
outpp7L13(11)<=outpp7L17(11);
outpp8L13(11)<=outpp8L17(11);
outpp9L13(11)<=outpp9L17(11);
outpp10L13(11)<=outpp10L17(11);
outpp11L13(11)<=outpp11L17(11);
outpp12L13(11)<=outpp12L17(11);
outpp0L13(12)<=outpp0L17(12);
outpp1L13(12)<=outpp1L17(12);
outpp2L13(12)<=outpp2L17(12);
outpp3L13(12)<=outpp3L17(12);
outpp4L13(12)<=outpp4L17(12);
outpp5L13(12)<=outpp5L17(12);
outpp6L13(12)<=outpp6L17(12);
outpp7L13(12)<=outpp7L17(12);
outpp8L13(12)<=outpp8L17(12);
outpp9L13(12)<=outpp9L17(12);
outpp10L13(12)<=outpp10L17(12);
outpp11L13(12)<=outpp11L17(12);
outpp12L13(12)<=outpp12L17(12);
outpp0L13(13)<=outpp0L17(13);
outpp1L13(13)<=outpp1L17(13);
outpp2L13(13)<=outpp2L17(13);
outpp3L13(13)<=outpp3L17(13);
outpp4L13(13)<=outpp4L17(13);
outpp5L13(13)<=outpp5L17(13);
outpp6L13(13)<=outpp6L17(13);
outpp7L13(13)<=outpp7L17(13);
outpp8L13(13)<=outpp8L17(13);
outpp9L13(13)<=outpp9L17(13);
outpp10L13(13)<=outpp10L17(13);
outpp11L13(13)<=outpp11L17(13);
outpp12L13(13)<=outpp12L17(13);
outpp0L13(14)<=outpp0L17(14);
outpp1L13(14)<=outpp1L17(14);
outpp2L13(14)<=outpp2L17(14);
outpp3L13(14)<=outpp3L17(14);
outpp4L13(14)<=outpp4L17(14);
outpp5L13(14)<=outpp5L17(14);
outpp6L13(14)<=outpp6L17(14);
outpp7L13(14)<=outpp7L17(14);
outpp8L13(14)<=outpp8L17(14);
outpp9L13(14)<=outpp9L17(14);
outpp10L13(14)<=outpp10L17(14);
outpp11L13(14)<=outpp11L17(14);
outpp12L13(14)<=outpp12L17(14);
outpp0L13(15)<=outpp0L17(15);
outpp1L13(15)<=outpp1L17(15);
outpp2L13(15)<=outpp2L17(15);
outpp3L13(15)<=outpp3L17(15);
outpp4L13(15)<=outpp4L17(15);
outpp5L13(15)<=outpp5L17(15);
outpp6L13(15)<=outpp6L17(15);
outpp7L13(15)<=outpp7L17(15);
outpp8L13(15)<=outpp8L17(15);
outpp9L13(15)<=outpp9L17(15);
outpp10L13(15)<=outpp10L17(15);
outpp11L13(15)<=outpp11L17(15);
outpp12L13(15)<=outpp12L17(15);
outpp0L13(16)<=outpp0L17(16);
outpp1L13(16)<=outpp1L17(16);
outpp2L13(16)<=outpp2L17(16);
outpp3L13(16)<=outpp3L17(16);
outpp4L13(16)<=outpp4L17(16);
outpp5L13(16)<=outpp5L17(16);
outpp6L13(16)<=outpp6L17(16);
outpp7L13(16)<=outpp7L17(16);
outpp8L13(16)<=outpp8L17(16);
outpp9L13(16)<=outpp9L17(16);
outpp10L13(16)<=outpp10L17(16);
outpp11L13(16)<=outpp11L17(16);
outpp12L13(16)<=outpp12L17(16);
outpp0L13(17)<=outpp0L17(17);
outpp1L13(17)<=outpp1L17(17);
outpp2L13(17)<=outpp2L17(17);
outpp3L13(17)<=outpp3L17(17);
outpp4L13(17)<=outpp4L17(17);
outpp5L13(17)<=outpp5L17(17);
outpp6L13(17)<=outpp6L17(17);
outpp7L13(17)<=outpp7L17(17);
outpp8L13(17)<=outpp8L17(17);
outpp9L13(17)<=outpp9L17(17);
outpp10L13(17)<=outpp10L17(17);
outpp11L13(17)<=outpp11L17(17);
outpp12L13(17)<=outpp12L17(17);
outpp0L13(18)<=outpp0L17(18);
outpp1L13(18)<=outpp1L17(18);
outpp2L13(18)<=outpp2L17(18);
outpp3L13(18)<=outpp3L17(18);
outpp4L13(18)<=outpp4L17(18);
outpp5L13(18)<=outpp5L17(18);
outpp6L13(18)<=outpp6L17(18);
outpp7L13(18)<=outpp7L17(18);
outpp8L13(18)<=outpp8L17(18);
outpp9L13(18)<=outpp9L17(18);
outpp10L13(18)<=outpp10L17(18);
outpp11L13(18)<=outpp11L17(18);
outpp12L13(18)<=outpp12L17(18);
outpp0L13(19)<=outpp0L17(19);
outpp1L13(19)<=outpp1L17(19);
outpp2L13(19)<=outpp2L17(19);
outpp3L13(19)<=outpp3L17(19);
outpp4L13(19)<=outpp4L17(19);
outpp5L13(19)<=outpp5L17(19);
outpp6L13(19)<=outpp6L17(19);
outpp7L13(19)<=outpp7L17(19);
outpp8L13(19)<=outpp8L17(19);
outpp9L13(19)<=outpp9L17(19);
outpp10L13(19)<=outpp10L17(19);
outpp11L13(19)<=outpp11L17(19);
outpp12L13(19)<=outpp12L17(19);
outpp0L13(20)<=outpp0L17(20);
outpp1L13(20)<=outpp1L17(20);
outpp2L13(20)<=outpp2L17(20);
outpp3L13(20)<=outpp3L17(20);
outpp4L13(20)<=outpp4L17(20);
outpp5L13(20)<=outpp5L17(20);
outpp6L13(20)<=outpp6L17(20);
outpp7L13(20)<=outpp7L17(20);
outpp8L13(20)<=outpp8L17(20);
outpp9L13(20)<=outpp9L17(20);
outpp10L13(20)<=outpp10L17(20);
outpp11L13(20)<=outpp11L17(20);
outpp12L13(20)<=outpp12L17(20);
outpp0L13(21)<=outpp0L17(21);
outpp1L13(21)<=outpp1L17(21);
outpp2L13(21)<=outpp2L17(21);
outpp3L13(21)<=outpp3L17(21);
outpp4L13(21)<=outpp4L17(21);
outpp5L13(21)<=outpp5L17(21);
outpp6L13(21)<=outpp6L17(21);
outpp7L13(21)<=outpp7L17(21);
outpp8L13(21)<=outpp8L17(21);
outpp9L13(21)<=outpp9L17(21);
outpp10L13(21)<=outpp10L17(21);
outpp11L13(21)<=outpp11L17(21);
outpp12L13(21)<=outpp12L17(21);
outpp0L13(22)<=outpp0L17(22);
outpp1L13(22)<=outpp1L17(22);
outpp2L13(22)<=outpp2L17(22);
outpp3L13(22)<=outpp3L17(22);
outpp4L13(22)<=outpp4L17(22);
outpp5L13(22)<=outpp5L17(22);
outpp6L13(22)<=outpp6L17(22);
outpp7L13(22)<=outpp7L17(22);
outpp8L13(22)<=outpp8L17(22);
outpp9L13(22)<=outpp9L17(22);
outpp10L13(22)<=outpp10L17(22);
outpp11L13(22)<=outpp11L17(22);
outpp12L13(22)<=outpp12L17(22);
outpp0L13(23)<=outpp0L17(23);
outpp1L13(23)<=outpp1L17(23);
outpp2L13(23)<=outpp2L17(23);
outpp3L13(23)<=outpp3L17(23);
outpp4L13(23)<=outpp4L17(23);
outpp5L13(23)<=outpp5L17(23);
outpp6L13(23)<=outpp6L17(23);
outpp7L13(23)<=outpp7L17(23);
outpp8L13(23)<=outpp8L17(23);
outpp9L13(23)<=outpp9L17(23);
outpp10L13(23)<=outpp10L17(23);
outpp11L13(23)<=outpp11L17(23);
outpp12L13(23)<=outpp12L17(23);
HA0L17: HA port map( A=>outpp0L17(24), B=>outpp1L17(24), S=>outpp0L13(24) ,cout=>outpp0L13(25));
outpp1L13(24)<=outpp2L17(24);
outpp2L13(24)<=outpp3L17(24);
outpp3L13(24)<=outpp4L17(24);
outpp4L13(24)<=outpp5L17(24);
outpp5L13(24)<=outpp6L17(24);
outpp6L13(24)<=outpp7L17(24);
outpp7L13(24)<=outpp8L17(24);
outpp8L13(24)<=outpp9L17(24);
outpp9L13(24)<=outpp10L17(24);
outpp10L13(24)<=outpp11L17(24);
outpp11L13(24)<=outpp12L17(24);
outpp12L13(24)<=outpp13L17(24);
HA1L17: HA port map( A=>outpp0L17(25), B=>outpp1L17(25), S=>outpp1L13(25) ,cout=>outpp0L13(26));
outpp2L13(25)<=outpp2L17(25);
outpp3L13(25)<=outpp3L17(25);
outpp4L13(25)<=outpp4L17(25);
outpp5L13(25)<=outpp5L17(25);
outpp6L13(25)<=outpp6L17(25);
outpp7L13(25)<=outpp7L17(25);
outpp8L13(25)<=outpp8L17(25);
outpp9L13(25)<=outpp9L17(25);
outpp10L13(25)<=outpp10L17(25);
outpp11L13(25)<=outpp11L17(25);
outpp12L13(25)<=outpp12L17(25);
HA2L17: HA port map( A=>outpp0L17(26), B=>outpp1L17(26), S=>outpp1L13(26) ,cout=>outpp0L13(27));
FA0L17: FA port map(A=>outpp2L17(26), B=>outpp3L17(26), cin=>outpp4L17(26), S=>outpp2L13(26) ,cout=>outpp1L13(27));
outpp3L13(26)<=outpp5L17(26);
outpp4L13(26)<=outpp6L17(26);
outpp5L13(26)<=outpp7L17(26);
outpp6L13(26)<=outpp8L17(26);
outpp7L13(26)<=outpp9L17(26);
outpp8L13(26)<=outpp10L17(26);
outpp9L13(26)<=outpp11L17(26);
outpp10L13(26)<=outpp12L17(26);
outpp11L13(26)<=outpp13L17(26);
outpp12L13(26)<=outpp14L17(26);
HA3L17: HA port map( A=>outpp0L17(27), B=>outpp1L17(27), S=>outpp2L13(27) ,cout=>outpp0L13(28));
FA1L17: FA port map(A=>outpp2L17(27), B=>outpp3L17(27), cin=>outpp4L17(27), S=>outpp3L13(27) ,cout=>outpp1L13(28));
outpp4L13(27)<=outpp5L17(27);
outpp5L13(27)<=outpp6L17(27);
outpp6L13(27)<=outpp7L17(27);
outpp7L13(27)<=outpp8L17(27);
outpp8L13(27)<=outpp9L17(27);
outpp9L13(27)<=outpp10L17(27);
outpp10L13(27)<=outpp11L17(27);
outpp11L13(27)<=outpp12L17(27);
outpp12L13(27)<=outpp13L17(27);
HA4L17: HA port map( A=>outpp0L17(28), B=>outpp1L17(28), S=>outpp2L13(28) ,cout=>outpp0L13(29));
FA2L17: FA port map(A=>outpp2L17(28), B=>outpp3L17(28), cin=>outpp4L17(28), S=>outpp3L13(28) ,cout=>outpp1L13(29));
FA3L17: FA port map(A=>outpp5L17(28), B=>outpp6L17(28), cin=>outpp7L17(28), S=>outpp4L13(28) ,cout=>outpp2L13(29));
outpp5L13(28)<=outpp8L17(28);
outpp6L13(28)<=outpp9L17(28);
outpp7L13(28)<=outpp10L17(28);
outpp8L13(28)<=outpp11L17(28);
outpp9L13(28)<=outpp12L17(28);
outpp10L13(28)<=outpp13L17(28);
outpp11L13(28)<=outpp14L17(28);
outpp12L13(28)<=outpp15L17(28);
HA5L17: HA port map( A=>outpp0L17(29), B=>outpp1L17(29), S=>outpp3L13(29) ,cout=>outpp0L13(30));
FA4L17: FA port map(A=>outpp2L17(29), B=>outpp3L17(29), cin=>outpp4L17(29), S=>outpp4L13(29) ,cout=>outpp1L13(30));
FA5L17: FA port map(A=>outpp5L17(29), B=>outpp6L17(29), cin=>outpp7L17(29), S=>outpp5L13(29) ,cout=>outpp2L13(30));
outpp6L13(29)<=outpp8L17(29);
outpp7L13(29)<=outpp9L17(29);
outpp8L13(29)<=outpp10L17(29);
outpp9L13(29)<=outpp11L17(29);
outpp10L13(29)<=outpp12L17(29);
outpp11L13(29)<=outpp13L17(29);
outpp12L13(29)<=outpp14L17(29);
HA6L17: HA port map( A=>outpp0L17(30), B=>outpp1L17(30), S=>outpp3L13(30) ,cout=>outpp0L13(31));
FA6L17: FA port map(A=>outpp2L17(30), B=>outpp3L17(30), cin=>outpp4L17(30), S=>outpp4L13(30) ,cout=>outpp1L13(31));
FA7L17: FA port map(A=>outpp5L17(30), B=>outpp6L17(30), cin=>outpp7L17(30), S=>outpp5L13(30) ,cout=>outpp2L13(31));
FA8L17: FA port map(A=>outpp8L17(30), B=>outpp9L17(30), cin=>outpp10L17(30), S=>outpp6L13(30) ,cout=>outpp3L13(31));
outpp7L13(30)<=outpp11L17(30);
outpp8L13(30)<=outpp12L17(30);
outpp9L13(30)<=outpp13L17(30);
outpp10L13(30)<=outpp14L17(30);
outpp11L13(30)<=outpp15L17(30);
outpp12L13(30)<=outpp16L17(30);
HA7L17: HA port map( A=>outpp0L17(31), B=>outpp1L17(31), S=>outpp4L13(31) ,cout=>outpp0L13(32));
FA9L17: FA port map(A=>outpp2L17(31), B=>outpp3L17(31), cin=>outpp4L17(31), S=>outpp5L13(31) ,cout=>outpp1L13(32));
FA10L17: FA port map(A=>outpp5L17(31), B=>outpp6L17(31), cin=>outpp7L17(31), S=>outpp6L13(31) ,cout=>outpp2L13(32));
FA11L17: FA port map(A=>outpp8L17(31), B=>outpp9L17(31), cin=>outpp10L17(31), S=>outpp7L13(31) ,cout=>outpp3L13(32));
outpp8L13(31)<=outpp11L17(31);
outpp9L13(31)<=outpp12L17(31);
outpp10L13(31)<=outpp13L17(31);
outpp11L13(31)<=outpp14L17(31);
outpp12L13(31)<=outpp15L17(31);
FA12L17: FA port map(A=>outpp0L17(32), B=>outpp1L17(32), cin=>outpp2L17(32), S=>outpp4L13(32) ,cout=>outpp0L13(33));
FA13L17: FA port map(A=>outpp3L17(32), B=>outpp4L17(32), cin=>outpp5L17(32), S=>outpp5L13(32) ,cout=>outpp1L13(33));
FA14L17: FA port map(A=>outpp6L17(32), B=>outpp7L17(32), cin=>outpp8L17(32), S=>outpp6L13(32) ,cout=>outpp2L13(33));
FA15L17: FA port map(A=>outpp9L17(32), B=>outpp10L17(32), cin=>outpp11L17(32), S=>outpp7L13(32) ,cout=>outpp3L13(33));
outpp8L13(32)<=outpp12L17(32);
outpp9L13(32)<=outpp13L17(32);
outpp10L13(32)<=outpp14L17(32);
outpp11L13(32)<=outpp15L17(32);
outpp12L13(32)<=outpp16L17(32);
FA16L17: FA port map(A=>outpp0L17(33), B=>outpp1L17(33), cin=>outpp2L17(33), S=>outpp4L13(33) ,cout=>outpp0L13(34));
FA17L17: FA port map(A=>outpp3L17(33), B=>outpp4L17(33), cin=>outpp5L17(33), S=>outpp5L13(33) ,cout=>outpp1L13(34));
FA18L17: FA port map(A=>outpp6L17(33), B=>outpp7L17(33), cin=>outpp8L17(33), S=>outpp6L13(33) ,cout=>outpp2L13(34));
FA19L17: FA port map(A=>outpp9L17(33), B=>outpp10L17(33), cin=>outpp11L17(33), S=>outpp7L13(33) ,cout=>outpp3L13(34));
outpp8L13(33)<=outpp12L17(33);
outpp9L13(33)<=outpp13L17(33);
outpp10L13(33)<=outpp14L17(33);
outpp11L13(33)<=outpp15L17(33);
outpp12L13(33)<=outpp16L17(33);
FA20L17: FA port map(A=>outpp0L17(34), B=>outpp1L17(34), cin=>outpp2L17(34), S=>outpp4L13(34) ,cout=>outpp0L13(35));
FA21L17: FA port map(A=>outpp3L17(34), B=>outpp4L17(34), cin=>outpp5L17(34), S=>outpp5L13(34) ,cout=>outpp1L13(35));
FA22L17: FA port map(A=>outpp6L17(34), B=>outpp7L17(34), cin=>outpp8L17(34), S=>outpp6L13(34) ,cout=>outpp2L13(35));
FA23L17: FA port map(A=>outpp9L17(34), B=>outpp10L17(34), cin=>outpp11L17(34), S=>outpp7L13(34) ,cout=>outpp3L13(35));
outpp8L13(34)<=outpp12L17(34);
outpp9L13(34)<=outpp13L17(34);
outpp10L13(34)<=outpp14L17(34);
outpp11L13(34)<=outpp15L17(34);
outpp12L13(34)<=outpp16L17(34);
FA24L17: FA port map(A=>outpp0L17(35), B=>outpp1L17(35), cin=>outpp2L17(35), S=>outpp4L13(35) ,cout=>outpp0L13(36));
FA25L17: FA port map(A=>outpp3L17(35), B=>outpp4L17(35), cin=>outpp5L17(35), S=>outpp5L13(35) ,cout=>outpp1L13(36));
FA26L17: FA port map(A=>outpp6L17(35), B=>outpp7L17(35), cin=>outpp8L17(35), S=>outpp6L13(35) ,cout=>outpp2L13(36));
FA27L17: FA port map(A=>outpp9L17(35), B=>outpp10L17(35), cin=>outpp11L17(35), S=>outpp7L13(35) ,cout=>outpp3L13(36));
outpp8L13(35)<=outpp12L17(35);
outpp9L13(35)<=outpp13L17(35);
outpp10L13(35)<=outpp14L17(35);
outpp11L13(35)<=outpp15L17(35);
outpp12L13(35)<=outpp16L17(35);
HA8L17: HA port map( A=>outpp1L17(36), B=>outpp2L17(36), S=>outpp4L13(36) ,cout=>outpp0L13(37));
FA28L17: FA port map(A=>outpp3L17(36), B=>outpp4L17(36), cin=>outpp5L17(36), S=>outpp5L13(36) ,cout=>outpp1L13(37));
FA29L17: FA port map(A=>outpp6L17(36), B=>outpp7L17(36), cin=>outpp8L17(36), S=>outpp6L13(36) ,cout=>outpp2L13(37));
FA30L17: FA port map(A=>outpp9L17(36), B=>outpp10L17(36), cin=>outpp11L17(36), S=>outpp7L13(36) ,cout=>outpp3L13(37));
outpp8L13(36)<=outpp12L17(36);
outpp9L13(36)<=outpp13L17(36);
outpp10L13(36)<=outpp14L17(36);
outpp11L13(36)<=outpp15L17(36);
outpp12L13(36)<=outpp16L17(36);
FA31L17: FA port map(A=>outpp2L17(37), B=>outpp3L17(37), cin=>outpp4L17(37), S=>outpp4L13(37) ,cout=>outpp0L13(38));
FA32L17: FA port map(A=>outpp5L17(37), B=>outpp6L17(37), cin=>outpp7L17(37), S=>outpp5L13(37) ,cout=>outpp1L13(38));
FA33L17: FA port map(A=>outpp8L17(37), B=>outpp9L17(37), cin=>outpp10L17(37), S=>outpp6L13(37) ,cout=>outpp2L13(38));
outpp7L13(37)<=outpp11L17(37);
outpp8L13(37)<=outpp12L17(37);
outpp9L13(37)<=outpp13L17(37);
outpp10L13(37)<=outpp14L17(37);
outpp11L13(37)<=outpp15L17(37);
outpp12L13(37)<=outpp16L17(37);
HA9L17: HA port map( A=>outpp2L17(38), B=>outpp3L17(38), S=>outpp3L13(38) ,cout=>outpp0L13(39));
FA34L17: FA port map(A=>outpp4L17(38), B=>outpp5L17(38), cin=>outpp6L17(38), S=>outpp4L13(38) ,cout=>outpp1L13(39));
FA35L17: FA port map(A=>outpp7L17(38), B=>outpp8L17(38), cin=>outpp9L17(38), S=>outpp5L13(38) ,cout=>outpp2L13(39));
outpp6L13(38)<=outpp10L17(38);
outpp7L13(38)<=outpp11L17(38);
outpp8L13(38)<=outpp12L17(38);
outpp9L13(38)<=outpp13L17(38);
outpp10L13(38)<=outpp14L17(38);
outpp11L13(38)<=outpp15L17(38);
outpp12L13(38)<=outpp16L17(38);
FA36L17: FA port map(A=>outpp3L17(39), B=>outpp4L17(39), cin=>outpp5L17(39), S=>outpp3L13(39) ,cout=>outpp0L13(40));
FA37L17: FA port map(A=>outpp6L17(39), B=>outpp7L17(39), cin=>outpp8L17(39), S=>outpp4L13(39) ,cout=>outpp1L13(40));
outpp5L13(39)<=outpp9L17(39);
outpp6L13(39)<=outpp10L17(39);
outpp7L13(39)<=outpp11L17(39);
outpp8L13(39)<=outpp12L17(39);
outpp9L13(39)<=outpp13L17(39);
outpp10L13(39)<=outpp14L17(39);
outpp11L13(39)<=outpp15L17(39);
outpp12L13(39)<=outpp16L17(39);
HA10L17: HA port map( A=>outpp3L17(40), B=>outpp4L17(40), S=>outpp2L13(40) ,cout=>outpp0L13(41));
FA38L17: FA port map(A=>outpp5L17(40), B=>outpp6L17(40), cin=>outpp7L17(40), S=>outpp3L13(40) ,cout=>outpp1L13(41));
outpp4L13(40)<=outpp8L17(40);
outpp5L13(40)<=outpp9L17(40);
outpp6L13(40)<=outpp10L17(40);
outpp7L13(40)<=outpp11L17(40);
outpp8L13(40)<=outpp12L17(40);
outpp9L13(40)<=outpp13L17(40);
outpp10L13(40)<=outpp14L17(40);
outpp11L13(40)<=outpp15L17(40);
outpp12L13(40)<=outpp16L17(40);
FA39L17: FA port map(A=>outpp4L17(41), B=>outpp5L17(41), cin=>outpp6L17(41), S=>outpp2L13(41) ,cout=>outpp0L13(42));
outpp3L13(41)<=outpp7L17(41);
outpp4L13(41)<=outpp8L17(41);
outpp5L13(41)<=outpp9L17(41);
outpp6L13(41)<=outpp10L17(41);
outpp7L13(41)<=outpp11L17(41);
outpp8L13(41)<=outpp12L17(41);
outpp9L13(41)<=outpp13L17(41);
outpp10L13(41)<=outpp14L17(41);
outpp11L13(41)<=outpp15L17(41);
outpp12L13(41)<=outpp16L17(41);
HA11L17: HA port map( A=>outpp4L17(42), B=>outpp5L17(42), S=>outpp1L13(42) ,cout=>outpp0L13(43));
outpp2L13(42)<=outpp6L17(42);
outpp3L13(42)<=outpp7L17(42);
outpp4L13(42)<=outpp8L17(42);
outpp5L13(42)<=outpp9L17(42);
outpp6L13(42)<=outpp10L17(42);
outpp7L13(42)<=outpp11L17(42);
outpp8L13(42)<=outpp12L17(42);
outpp9L13(42)<=outpp13L17(42);
outpp10L13(42)<=outpp14L17(42);
outpp11L13(42)<=outpp15L17(42);
outpp12L13(42)<=outpp16L17(42);
outpp1L13(43)<=outpp5L17(43);
outpp2L13(43)<=outpp6L17(43);
outpp3L13(43)<=outpp7L17(43);
outpp4L13(43)<=outpp8L17(43);
outpp5L13(43)<=outpp9L17(43);
outpp6L13(43)<=outpp10L17(43);
outpp7L13(43)<=outpp11L17(43);
outpp8L13(43)<=outpp12L17(43);
outpp9L13(43)<=outpp13L17(43);
outpp10L13(43)<=outpp14L17(43);
outpp11L13(43)<=outpp15L17(43);
outpp12L13(43)<=outpp16L17(43);
outpp0L13(44)<=outpp5L17(44);
outpp1L13(44)<=outpp6L17(44);
outpp2L13(44)<=outpp7L17(44);
outpp3L13(44)<=outpp8L17(44);
outpp4L13(44)<=outpp9L17(44);
outpp5L13(44)<=outpp10L17(44);
outpp6L13(44)<=outpp11L17(44);
outpp7L13(44)<=outpp12L17(44);
outpp8L13(44)<=outpp13L17(44);
outpp9L13(44)<=outpp14L17(44);
outpp10L13(44)<=outpp15L17(44);
outpp11L13(44)<=outpp16L17(44);
outpp0L13(45)<=outpp6L17(45);
outpp1L13(45)<=outpp7L17(45);
outpp2L13(45)<=outpp8L17(45);
outpp3L13(45)<=outpp9L17(45);
outpp4L13(45)<=outpp10L17(45);
outpp5L13(45)<=outpp11L17(45);
outpp6L13(45)<=outpp12L17(45);
outpp7L13(45)<=outpp13L17(45);
outpp8L13(45)<=outpp14L17(45);
outpp9L13(45)<=outpp15L17(45);
outpp10L13(45)<=outpp16L17(45);
outpp0L13(46)<=outpp6L17(46);
outpp1L13(46)<=outpp7L17(46);
outpp2L13(46)<=outpp8L17(46);
outpp3L13(46)<=outpp9L17(46);
outpp4L13(46)<=outpp10L17(46);
outpp5L13(46)<=outpp11L17(46);
outpp6L13(46)<=outpp12L17(46);
outpp7L13(46)<=outpp13L17(46);
outpp8L13(46)<=outpp14L17(46);
outpp9L13(46)<=outpp15L17(46);
outpp10L13(46)<=outpp16L17(46);
outpp0L13(47)<=outpp7L17(47);
outpp1L13(47)<=outpp8L17(47);
outpp2L13(47)<=outpp9L17(47);
outpp3L13(47)<=outpp10L17(47);
outpp4L13(47)<=outpp11L17(47);
outpp5L13(47)<=outpp12L17(47);
outpp6L13(47)<=outpp13L17(47);
outpp7L13(47)<=outpp14L17(47);
outpp8L13(47)<=outpp15L17(47);
outpp9L13(47)<=outpp16L17(47);
outpp0L13(48)<=outpp7L17(48);
outpp1L13(48)<=outpp8L17(48);
outpp2L13(48)<=outpp9L17(48);
outpp3L13(48)<=outpp10L17(48);
outpp4L13(48)<=outpp11L17(48);
outpp5L13(48)<=outpp12L17(48);
outpp6L13(48)<=outpp13L17(48);
outpp7L13(48)<=outpp14L17(48);
outpp8L13(48)<=outpp15L17(48);
outpp9L13(48)<=outpp16L17(48);
outpp0L13(49)<=outpp8L17(49);
outpp1L13(49)<=outpp9L17(49);
outpp2L13(49)<=outpp10L17(49);
outpp3L13(49)<=outpp11L17(49);
outpp4L13(49)<=outpp12L17(49);
outpp5L13(49)<=outpp13L17(49);
outpp6L13(49)<=outpp14L17(49);
outpp7L13(49)<=outpp15L17(49);
outpp8L13(49)<=outpp16L17(49);
outpp0L13(50)<=outpp8L17(50);
outpp1L13(50)<=outpp9L17(50);
outpp2L13(50)<=outpp10L17(50);
outpp3L13(50)<=outpp11L17(50);
outpp4L13(50)<=outpp12L17(50);
outpp5L13(50)<=outpp13L17(50);
outpp6L13(50)<=outpp14L17(50);
outpp7L13(50)<=outpp15L17(50);
outpp8L13(50)<=outpp16L17(50);
outpp0L13(51)<=outpp9L17(51);
outpp1L13(51)<=outpp10L17(51);
outpp2L13(51)<=outpp11L17(51);
outpp3L13(51)<=outpp12L17(51);
outpp4L13(51)<=outpp13L17(51);
outpp5L13(51)<=outpp14L17(51);
outpp6L13(51)<=outpp15L17(51);
outpp7L13(51)<=outpp16L17(51);
outpp0L13(52)<=outpp9L17(52);
outpp1L13(52)<=outpp10L17(52);
outpp2L13(52)<=outpp11L17(52);
outpp3L13(52)<=outpp12L17(52);
outpp4L13(52)<=outpp13L17(52);
outpp5L13(52)<=outpp14L17(52);
outpp6L13(52)<=outpp15L17(52);
outpp7L13(52)<=outpp16L17(52);
outpp0L13(53)<=outpp10L17(53);
outpp1L13(53)<=outpp11L17(53);
outpp2L13(53)<=outpp12L17(53);
outpp3L13(53)<=outpp13L17(53);
outpp4L13(53)<=outpp14L17(53);
outpp5L13(53)<=outpp15L17(53);
outpp6L13(53)<=outpp16L17(53);
outpp0L13(54)<=outpp10L17(54);
outpp1L13(54)<=outpp11L17(54);
outpp2L13(54)<=outpp12L17(54);
outpp3L13(54)<=outpp13L17(54);
outpp4L13(54)<=outpp14L17(54);
outpp5L13(54)<=outpp15L17(54);
outpp6L13(54)<=outpp16L17(54);
outpp0L13(55)<=outpp11L17(55);
outpp1L13(55)<=outpp12L17(55);
outpp2L13(55)<=outpp13L17(55);
outpp3L13(55)<=outpp14L17(55);
outpp4L13(55)<=outpp15L17(55);
outpp5L13(55)<=outpp16L17(55);
outpp0L13(56)<=outpp11L17(56);
outpp1L13(56)<=outpp12L17(56);
outpp2L13(56)<=outpp13L17(56);
outpp3L13(56)<=outpp14L17(56);
outpp4L13(56)<=outpp15L17(56);
outpp5L13(56)<=outpp16L17(56);
outpp0L13(57)<=outpp12L17(57);
outpp1L13(57)<=outpp13L17(57);
outpp2L13(57)<=outpp14L17(57);
outpp3L13(57)<=outpp15L17(57);
outpp4L13(57)<=outpp16L17(57);
outpp0L13(58)<=outpp12L17(58);
outpp1L13(58)<=outpp13L17(58);
outpp2L13(58)<=outpp14L17(58);
outpp3L13(58)<=outpp15L17(58);
outpp4L13(58)<=outpp16L17(58);
outpp0L13(59)<=outpp13L17(59);
outpp1L13(59)<=outpp14L17(59);
outpp2L13(59)<=outpp15L17(59);
outpp3L13(59)<=outpp16L17(59);
outpp0L13(60)<=outpp13L17(60);
outpp1L13(60)<=outpp14L17(60);
outpp2L13(60)<=outpp15L17(60);
outpp3L13(60)<=outpp16L17(60);
outpp0L13(61)<=outpp14L17(61);
outpp1L13(61)<=outpp15L17(61);
outpp2L13(61)<=outpp16L17(61);
outpp0L13(62)<=outpp14L17(62);
outpp1L13(62)<=outpp15L17(62);
outpp2L13(62)<=outpp16L17(62);
outpp0L13(63)<=outpp15L17(63);
outpp1L13(63)<=outpp16L17(63);
outpp0L9(0)<=outpp0L13(0);
outpp1L9(0)<=outpp1L13(0);
outpp2L9(0)<=outpp2L13(0);
outpp3L9(0)<=outpp3L13(0);
outpp4L9(0)<=outpp4L13(0);
outpp5L9(0)<=outpp5L13(0);
outpp6L9(0)<=outpp6L13(0);
outpp7L9(0)<=outpp7L13(0);
outpp8L9(0)<=outpp8L13(0);
outpp0L9(1)<=outpp0L13(1);
outpp1L9(1)<=outpp1L13(1);
outpp2L9(1)<=outpp2L13(1);
outpp3L9(1)<=outpp3L13(1);
outpp4L9(1)<=outpp4L13(1);
outpp5L9(1)<=outpp5L13(1);
outpp6L9(1)<=outpp6L13(1);
outpp7L9(1)<=outpp7L13(1);
outpp8L9(1)<=outpp8L13(1);
outpp0L9(2)<=outpp0L13(2);
outpp1L9(2)<=outpp1L13(2);
outpp2L9(2)<=outpp2L13(2);
outpp3L9(2)<=outpp3L13(2);
outpp4L9(2)<=outpp4L13(2);
outpp5L9(2)<=outpp5L13(2);
outpp6L9(2)<=outpp6L13(2);
outpp7L9(2)<=outpp7L13(2);
outpp8L9(2)<=outpp8L13(2);
outpp0L9(3)<=outpp0L13(3);
outpp1L9(3)<=outpp1L13(3);
outpp2L9(3)<=outpp2L13(3);
outpp3L9(3)<=outpp3L13(3);
outpp4L9(3)<=outpp4L13(3);
outpp5L9(3)<=outpp5L13(3);
outpp6L9(3)<=outpp6L13(3);
outpp7L9(3)<=outpp7L13(3);
outpp8L9(3)<=outpp8L13(3);
outpp0L9(4)<=outpp0L13(4);
outpp1L9(4)<=outpp1L13(4);
outpp2L9(4)<=outpp2L13(4);
outpp3L9(4)<=outpp3L13(4);
outpp4L9(4)<=outpp4L13(4);
outpp5L9(4)<=outpp5L13(4);
outpp6L9(4)<=outpp6L13(4);
outpp7L9(4)<=outpp7L13(4);
outpp8L9(4)<=outpp8L13(4);
outpp0L9(5)<=outpp0L13(5);
outpp1L9(5)<=outpp1L13(5);
outpp2L9(5)<=outpp2L13(5);
outpp3L9(5)<=outpp3L13(5);
outpp4L9(5)<=outpp4L13(5);
outpp5L9(5)<=outpp5L13(5);
outpp6L9(5)<=outpp6L13(5);
outpp7L9(5)<=outpp7L13(5);
outpp8L9(5)<=outpp8L13(5);
outpp0L9(6)<=outpp0L13(6);
outpp1L9(6)<=outpp1L13(6);
outpp2L9(6)<=outpp2L13(6);
outpp3L9(6)<=outpp3L13(6);
outpp4L9(6)<=outpp4L13(6);
outpp5L9(6)<=outpp5L13(6);
outpp6L9(6)<=outpp6L13(6);
outpp7L9(6)<=outpp7L13(6);
outpp8L9(6)<=outpp8L13(6);
outpp0L9(7)<=outpp0L13(7);
outpp1L9(7)<=outpp1L13(7);
outpp2L9(7)<=outpp2L13(7);
outpp3L9(7)<=outpp3L13(7);
outpp4L9(7)<=outpp4L13(7);
outpp5L9(7)<=outpp5L13(7);
outpp6L9(7)<=outpp6L13(7);
outpp7L9(7)<=outpp7L13(7);
outpp8L9(7)<=outpp8L13(7);
outpp0L9(8)<=outpp0L13(8);
outpp1L9(8)<=outpp1L13(8);
outpp2L9(8)<=outpp2L13(8);
outpp3L9(8)<=outpp3L13(8);
outpp4L9(8)<=outpp4L13(8);
outpp5L9(8)<=outpp5L13(8);
outpp6L9(8)<=outpp6L13(8);
outpp7L9(8)<=outpp7L13(8);
outpp8L9(8)<=outpp8L13(8);
outpp0L9(9)<=outpp0L13(9);
outpp1L9(9)<=outpp1L13(9);
outpp2L9(9)<=outpp2L13(9);
outpp3L9(9)<=outpp3L13(9);
outpp4L9(9)<=outpp4L13(9);
outpp5L9(9)<=outpp5L13(9);
outpp6L9(9)<=outpp6L13(9);
outpp7L9(9)<=outpp7L13(9);
outpp8L9(9)<=outpp8L13(9);
outpp0L9(10)<=outpp0L13(10);
outpp1L9(10)<=outpp1L13(10);
outpp2L9(10)<=outpp2L13(10);
outpp3L9(10)<=outpp3L13(10);
outpp4L9(10)<=outpp4L13(10);
outpp5L9(10)<=outpp5L13(10);
outpp6L9(10)<=outpp6L13(10);
outpp7L9(10)<=outpp7L13(10);
outpp8L9(10)<=outpp8L13(10);
outpp0L9(11)<=outpp0L13(11);
outpp1L9(11)<=outpp1L13(11);
outpp2L9(11)<=outpp2L13(11);
outpp3L9(11)<=outpp3L13(11);
outpp4L9(11)<=outpp4L13(11);
outpp5L9(11)<=outpp5L13(11);
outpp6L9(11)<=outpp6L13(11);
outpp7L9(11)<=outpp7L13(11);
outpp8L9(11)<=outpp8L13(11);
outpp0L9(12)<=outpp0L13(12);
outpp1L9(12)<=outpp1L13(12);
outpp2L9(12)<=outpp2L13(12);
outpp3L9(12)<=outpp3L13(12);
outpp4L9(12)<=outpp4L13(12);
outpp5L9(12)<=outpp5L13(12);
outpp6L9(12)<=outpp6L13(12);
outpp7L9(12)<=outpp7L13(12);
outpp8L9(12)<=outpp8L13(12);
outpp0L9(13)<=outpp0L13(13);
outpp1L9(13)<=outpp1L13(13);
outpp2L9(13)<=outpp2L13(13);
outpp3L9(13)<=outpp3L13(13);
outpp4L9(13)<=outpp4L13(13);
outpp5L9(13)<=outpp5L13(13);
outpp6L9(13)<=outpp6L13(13);
outpp7L9(13)<=outpp7L13(13);
outpp8L9(13)<=outpp8L13(13);
outpp0L9(14)<=outpp0L13(14);
outpp1L9(14)<=outpp1L13(14);
outpp2L9(14)<=outpp2L13(14);
outpp3L9(14)<=outpp3L13(14);
outpp4L9(14)<=outpp4L13(14);
outpp5L9(14)<=outpp5L13(14);
outpp6L9(14)<=outpp6L13(14);
outpp7L9(14)<=outpp7L13(14);
outpp8L9(14)<=outpp8L13(14);
outpp0L9(15)<=outpp0L13(15);
outpp1L9(15)<=outpp1L13(15);
outpp2L9(15)<=outpp2L13(15);
outpp3L9(15)<=outpp3L13(15);
outpp4L9(15)<=outpp4L13(15);
outpp5L9(15)<=outpp5L13(15);
outpp6L9(15)<=outpp6L13(15);
outpp7L9(15)<=outpp7L13(15);
outpp8L9(15)<=outpp8L13(15);
HA12L13: HA port map( A=>outpp0L13(16), B=>outpp1L13(16), S=>outpp0L9(16) ,cout=>outpp0L9(17));
outpp1L9(16)<=outpp2L13(16);
outpp2L9(16)<=outpp3L13(16);
outpp3L9(16)<=outpp4L13(16);
outpp4L9(16)<=outpp5L13(16);
outpp5L9(16)<=outpp6L13(16);
outpp6L9(16)<=outpp7L13(16);
outpp7L9(16)<=outpp8L13(16);
outpp8L9(16)<=outpp9L13(16);
HA13L13: HA port map( A=>outpp0L13(17), B=>outpp1L13(17), S=>outpp1L9(17) ,cout=>outpp0L9(18));
outpp2L9(17)<=outpp2L13(17);
outpp3L9(17)<=outpp3L13(17);
outpp4L9(17)<=outpp4L13(17);
outpp5L9(17)<=outpp5L13(17);
outpp6L9(17)<=outpp6L13(17);
outpp7L9(17)<=outpp7L13(17);
outpp8L9(17)<=outpp8L13(17);
HA14L13: HA port map( A=>outpp0L13(18), B=>outpp1L13(18), S=>outpp1L9(18) ,cout=>outpp0L9(19));
FA40L13: FA port map(A=>outpp2L13(18), B=>outpp3L13(18), cin=>outpp4L13(18), S=>outpp2L9(18) ,cout=>outpp1L9(19));
outpp3L9(18)<=outpp5L13(18);
outpp4L9(18)<=outpp6L13(18);
outpp5L9(18)<=outpp7L13(18);
outpp6L9(18)<=outpp8L13(18);
outpp7L9(18)<=outpp9L13(18);
outpp8L9(18)<=outpp10L13(18);
HA15L13: HA port map( A=>outpp0L13(19), B=>outpp1L13(19), S=>outpp2L9(19) ,cout=>outpp0L9(20));
FA41L13: FA port map(A=>outpp2L13(19), B=>outpp3L13(19), cin=>outpp4L13(19), S=>outpp3L9(19) ,cout=>outpp1L9(20));
outpp4L9(19)<=outpp5L13(19);
outpp5L9(19)<=outpp6L13(19);
outpp6L9(19)<=outpp7L13(19);
outpp7L9(19)<=outpp8L13(19);
outpp8L9(19)<=outpp9L13(19);
HA16L13: HA port map( A=>outpp0L13(20), B=>outpp1L13(20), S=>outpp2L9(20) ,cout=>outpp0L9(21));
FA42L13: FA port map(A=>outpp2L13(20), B=>outpp3L13(20), cin=>outpp4L13(20), S=>outpp3L9(20) ,cout=>outpp1L9(21));
FA43L13: FA port map(A=>outpp5L13(20), B=>outpp6L13(20), cin=>outpp7L13(20), S=>outpp4L9(20) ,cout=>outpp2L9(21));
outpp5L9(20)<=outpp8L13(20);
outpp6L9(20)<=outpp9L13(20);
outpp7L9(20)<=outpp10L13(20);
outpp8L9(20)<=outpp11L13(20);
HA17L13: HA port map( A=>outpp0L13(21), B=>outpp1L13(21), S=>outpp3L9(21) ,cout=>outpp0L9(22));
FA44L13: FA port map(A=>outpp2L13(21), B=>outpp3L13(21), cin=>outpp4L13(21), S=>outpp4L9(21) ,cout=>outpp1L9(22));
FA45L13: FA port map(A=>outpp5L13(21), B=>outpp6L13(21), cin=>outpp7L13(21), S=>outpp5L9(21) ,cout=>outpp2L9(22));
outpp6L9(21)<=outpp8L13(21);
outpp7L9(21)<=outpp9L13(21);
outpp8L9(21)<=outpp10L13(21);
HA18L13: HA port map( A=>outpp0L13(22), B=>outpp1L13(22), S=>outpp3L9(22) ,cout=>outpp0L9(23));
FA46L13: FA port map(A=>outpp2L13(22), B=>outpp3L13(22), cin=>outpp4L13(22), S=>outpp4L9(22) ,cout=>outpp1L9(23));
FA47L13: FA port map(A=>outpp5L13(22), B=>outpp6L13(22), cin=>outpp7L13(22), S=>outpp5L9(22) ,cout=>outpp2L9(23));
FA48L13: FA port map(A=>outpp8L13(22), B=>outpp9L13(22), cin=>outpp10L13(22), S=>outpp6L9(22) ,cout=>outpp3L9(23));
outpp7L9(22)<=outpp11L13(22);
outpp8L9(22)<=outpp12L13(22);
HA19L13: HA port map( A=>outpp0L13(23), B=>outpp1L13(23), S=>outpp4L9(23) ,cout=>outpp0L9(24));
FA49L13: FA port map(A=>outpp2L13(23), B=>outpp3L13(23), cin=>outpp4L13(23), S=>outpp5L9(23) ,cout=>outpp1L9(24));
FA50L13: FA port map(A=>outpp5L13(23), B=>outpp6L13(23), cin=>outpp7L13(23), S=>outpp6L9(23) ,cout=>outpp2L9(24));
FA51L13: FA port map(A=>outpp8L13(23), B=>outpp9L13(23), cin=>outpp10L13(23), S=>outpp7L9(23) ,cout=>outpp3L9(24));
outpp8L9(23)<=outpp11L13(23);
FA52L13: FA port map(A=>outpp0L13(24), B=>outpp1L13(24), cin=>outpp2L13(24), S=>outpp4L9(24) ,cout=>outpp0L9(25));
FA53L13: FA port map(A=>outpp3L13(24), B=>outpp4L13(24), cin=>outpp5L13(24), S=>outpp5L9(24) ,cout=>outpp1L9(25));
FA54L13: FA port map(A=>outpp6L13(24), B=>outpp7L13(24), cin=>outpp8L13(24), S=>outpp6L9(24) ,cout=>outpp2L9(25));
FA55L13: FA port map(A=>outpp9L13(24), B=>outpp10L13(24), cin=>outpp11L13(24), S=>outpp7L9(24) ,cout=>outpp3L9(25));
outpp8L9(24)<=outpp12L13(24);
FA56L13: FA port map(A=>outpp0L13(25), B=>outpp1L13(25), cin=>outpp2L13(25), S=>outpp4L9(25) ,cout=>outpp0L9(26));
FA57L13: FA port map(A=>outpp3L13(25), B=>outpp4L13(25), cin=>outpp5L13(25), S=>outpp5L9(25) ,cout=>outpp1L9(26));
FA58L13: FA port map(A=>outpp6L13(25), B=>outpp7L13(25), cin=>outpp8L13(25), S=>outpp6L9(25) ,cout=>outpp2L9(26));
FA59L13: FA port map(A=>outpp9L13(25), B=>outpp10L13(25), cin=>outpp11L13(25), S=>outpp7L9(25) ,cout=>outpp3L9(26));
outpp8L9(25)<=outpp12L13(25);
FA60L13: FA port map(A=>outpp0L13(26), B=>outpp1L13(26), cin=>outpp2L13(26), S=>outpp4L9(26) ,cout=>outpp0L9(27));
FA61L13: FA port map(A=>outpp3L13(26), B=>outpp4L13(26), cin=>outpp5L13(26), S=>outpp5L9(26) ,cout=>outpp1L9(27));
FA62L13: FA port map(A=>outpp6L13(26), B=>outpp7L13(26), cin=>outpp8L13(26), S=>outpp6L9(26) ,cout=>outpp2L9(27));
FA63L13: FA port map(A=>outpp9L13(26), B=>outpp10L13(26), cin=>outpp11L13(26), S=>outpp7L9(26) ,cout=>outpp3L9(27));
outpp8L9(26)<=outpp12L13(26);
FA64L13: FA port map(A=>outpp0L13(27), B=>outpp1L13(27), cin=>outpp2L13(27), S=>outpp4L9(27) ,cout=>outpp0L9(28));
FA65L13: FA port map(A=>outpp3L13(27), B=>outpp4L13(27), cin=>outpp5L13(27), S=>outpp5L9(27) ,cout=>outpp1L9(28));
FA66L13: FA port map(A=>outpp6L13(27), B=>outpp7L13(27), cin=>outpp8L13(27), S=>outpp6L9(27) ,cout=>outpp2L9(28));
FA67L13: FA port map(A=>outpp9L13(27), B=>outpp10L13(27), cin=>outpp11L13(27), S=>outpp7L9(27) ,cout=>outpp3L9(28));
outpp8L9(27)<=outpp12L13(27);
FA68L13: FA port map(A=>outpp0L13(28), B=>outpp1L13(28), cin=>outpp2L13(28), S=>outpp4L9(28) ,cout=>outpp0L9(29));
FA69L13: FA port map(A=>outpp3L13(28), B=>outpp4L13(28), cin=>outpp5L13(28), S=>outpp5L9(28) ,cout=>outpp1L9(29));
FA70L13: FA port map(A=>outpp6L13(28), B=>outpp7L13(28), cin=>outpp8L13(28), S=>outpp6L9(28) ,cout=>outpp2L9(29));
FA71L13: FA port map(A=>outpp9L13(28), B=>outpp10L13(28), cin=>outpp11L13(28), S=>outpp7L9(28) ,cout=>outpp3L9(29));
outpp8L9(28)<=outpp12L13(28);
FA72L13: FA port map(A=>outpp0L13(29), B=>outpp1L13(29), cin=>outpp2L13(29), S=>outpp4L9(29) ,cout=>outpp0L9(30));
FA73L13: FA port map(A=>outpp3L13(29), B=>outpp4L13(29), cin=>outpp5L13(29), S=>outpp5L9(29) ,cout=>outpp1L9(30));
FA74L13: FA port map(A=>outpp6L13(29), B=>outpp7L13(29), cin=>outpp8L13(29), S=>outpp6L9(29) ,cout=>outpp2L9(30));
FA75L13: FA port map(A=>outpp9L13(29), B=>outpp10L13(29), cin=>outpp11L13(29), S=>outpp7L9(29) ,cout=>outpp3L9(30));
outpp8L9(29)<=outpp12L13(29);
FA76L13: FA port map(A=>outpp0L13(30), B=>outpp1L13(30), cin=>outpp2L13(30), S=>outpp4L9(30) ,cout=>outpp0L9(31));
FA77L13: FA port map(A=>outpp3L13(30), B=>outpp4L13(30), cin=>outpp5L13(30), S=>outpp5L9(30) ,cout=>outpp1L9(31));
FA78L13: FA port map(A=>outpp6L13(30), B=>outpp7L13(30), cin=>outpp8L13(30), S=>outpp6L9(30) ,cout=>outpp2L9(31));
FA79L13: FA port map(A=>outpp9L13(30), B=>outpp10L13(30), cin=>outpp11L13(30), S=>outpp7L9(30) ,cout=>outpp3L9(31));
outpp8L9(30)<=outpp12L13(30);
FA80L13: FA port map(A=>outpp0L13(31), B=>outpp1L13(31), cin=>outpp2L13(31), S=>outpp4L9(31) ,cout=>outpp0L9(32));
FA81L13: FA port map(A=>outpp3L13(31), B=>outpp4L13(31), cin=>outpp5L13(31), S=>outpp5L9(31) ,cout=>outpp1L9(32));
FA82L13: FA port map(A=>outpp6L13(31), B=>outpp7L13(31), cin=>outpp8L13(31), S=>outpp6L9(31) ,cout=>outpp2L9(32));
FA83L13: FA port map(A=>outpp9L13(31), B=>outpp10L13(31), cin=>outpp11L13(31), S=>outpp7L9(31) ,cout=>outpp3L9(32));
outpp8L9(31)<=outpp12L13(31);
FA84L13: FA port map(A=>outpp0L13(32), B=>outpp1L13(32), cin=>outpp2L13(32), S=>outpp4L9(32) ,cout=>outpp0L9(33));
FA85L13: FA port map(A=>outpp3L13(32), B=>outpp4L13(32), cin=>outpp5L13(32), S=>outpp5L9(32) ,cout=>outpp1L9(33));
FA86L13: FA port map(A=>outpp6L13(32), B=>outpp7L13(32), cin=>outpp8L13(32), S=>outpp6L9(32) ,cout=>outpp2L9(33));
FA87L13: FA port map(A=>outpp9L13(32), B=>outpp10L13(32), cin=>outpp11L13(32), S=>outpp7L9(32) ,cout=>outpp3L9(33));
outpp8L9(32)<=outpp12L13(32);
FA88L13: FA port map(A=>outpp0L13(33), B=>outpp1L13(33), cin=>outpp2L13(33), S=>outpp4L9(33) ,cout=>outpp0L9(34));
FA89L13: FA port map(A=>outpp3L13(33), B=>outpp4L13(33), cin=>outpp5L13(33), S=>outpp5L9(33) ,cout=>outpp1L9(34));
FA90L13: FA port map(A=>outpp6L13(33), B=>outpp7L13(33), cin=>outpp8L13(33), S=>outpp6L9(33) ,cout=>outpp2L9(34));
FA91L13: FA port map(A=>outpp9L13(33), B=>outpp10L13(33), cin=>outpp11L13(33), S=>outpp7L9(33) ,cout=>outpp3L9(34));
outpp8L9(33)<=outpp12L13(33);
FA92L13: FA port map(A=>outpp0L13(34), B=>outpp1L13(34), cin=>outpp2L13(34), S=>outpp4L9(34) ,cout=>outpp0L9(35));
FA93L13: FA port map(A=>outpp3L13(34), B=>outpp4L13(34), cin=>outpp5L13(34), S=>outpp5L9(34) ,cout=>outpp1L9(35));
FA94L13: FA port map(A=>outpp6L13(34), B=>outpp7L13(34), cin=>outpp8L13(34), S=>outpp6L9(34) ,cout=>outpp2L9(35));
FA95L13: FA port map(A=>outpp9L13(34), B=>outpp10L13(34), cin=>outpp11L13(34), S=>outpp7L9(34) ,cout=>outpp3L9(35));
outpp8L9(34)<=outpp12L13(34);
FA96L13: FA port map(A=>outpp0L13(35), B=>outpp1L13(35), cin=>outpp2L13(35), S=>outpp4L9(35) ,cout=>outpp0L9(36));
FA97L13: FA port map(A=>outpp3L13(35), B=>outpp4L13(35), cin=>outpp5L13(35), S=>outpp5L9(35) ,cout=>outpp1L9(36));
FA98L13: FA port map(A=>outpp6L13(35), B=>outpp7L13(35), cin=>outpp8L13(35), S=>outpp6L9(35) ,cout=>outpp2L9(36));
FA99L13: FA port map(A=>outpp9L13(35), B=>outpp10L13(35), cin=>outpp11L13(35), S=>outpp7L9(35) ,cout=>outpp3L9(36));
outpp8L9(35)<=outpp12L13(35);
FA100L13: FA port map(A=>outpp0L13(36), B=>outpp1L13(36), cin=>outpp2L13(36), S=>outpp4L9(36) ,cout=>outpp0L9(37));
FA101L13: FA port map(A=>outpp3L13(36), B=>outpp4L13(36), cin=>outpp5L13(36), S=>outpp5L9(36) ,cout=>outpp1L9(37));
FA102L13: FA port map(A=>outpp6L13(36), B=>outpp7L13(36), cin=>outpp8L13(36), S=>outpp6L9(36) ,cout=>outpp2L9(37));
FA103L13: FA port map(A=>outpp9L13(36), B=>outpp10L13(36), cin=>outpp11L13(36), S=>outpp7L9(36) ,cout=>outpp3L9(37));
outpp8L9(36)<=outpp12L13(36);
FA104L13: FA port map(A=>outpp0L13(37), B=>outpp1L13(37), cin=>outpp2L13(37), S=>outpp4L9(37) ,cout=>outpp0L9(38));
FA105L13: FA port map(A=>outpp3L13(37), B=>outpp4L13(37), cin=>outpp5L13(37), S=>outpp5L9(37) ,cout=>outpp1L9(38));
FA106L13: FA port map(A=>outpp6L13(37), B=>outpp7L13(37), cin=>outpp8L13(37), S=>outpp6L9(37) ,cout=>outpp2L9(38));
FA107L13: FA port map(A=>outpp9L13(37), B=>outpp10L13(37), cin=>outpp11L13(37), S=>outpp7L9(37) ,cout=>outpp3L9(38));
outpp8L9(37)<=outpp12L13(37);
FA108L13: FA port map(A=>outpp0L13(38), B=>outpp1L13(38), cin=>outpp2L13(38), S=>outpp4L9(38) ,cout=>outpp0L9(39));
FA109L13: FA port map(A=>outpp3L13(38), B=>outpp4L13(38), cin=>outpp5L13(38), S=>outpp5L9(38) ,cout=>outpp1L9(39));
FA110L13: FA port map(A=>outpp6L13(38), B=>outpp7L13(38), cin=>outpp8L13(38), S=>outpp6L9(38) ,cout=>outpp2L9(39));
FA111L13: FA port map(A=>outpp9L13(38), B=>outpp10L13(38), cin=>outpp11L13(38), S=>outpp7L9(38) ,cout=>outpp3L9(39));
outpp8L9(38)<=outpp12L13(38);
FA112L13: FA port map(A=>outpp0L13(39), B=>outpp1L13(39), cin=>outpp2L13(39), S=>outpp4L9(39) ,cout=>outpp0L9(40));
FA113L13: FA port map(A=>outpp3L13(39), B=>outpp4L13(39), cin=>outpp5L13(39), S=>outpp5L9(39) ,cout=>outpp1L9(40));
FA114L13: FA port map(A=>outpp6L13(39), B=>outpp7L13(39), cin=>outpp8L13(39), S=>outpp6L9(39) ,cout=>outpp2L9(40));
FA115L13: FA port map(A=>outpp9L13(39), B=>outpp10L13(39), cin=>outpp11L13(39), S=>outpp7L9(39) ,cout=>outpp3L9(40));
outpp8L9(39)<=outpp12L13(39);
FA116L13: FA port map(A=>outpp0L13(40), B=>outpp1L13(40), cin=>outpp2L13(40), S=>outpp4L9(40) ,cout=>outpp0L9(41));
FA117L13: FA port map(A=>outpp3L13(40), B=>outpp4L13(40), cin=>outpp5L13(40), S=>outpp5L9(40) ,cout=>outpp1L9(41));
FA118L13: FA port map(A=>outpp6L13(40), B=>outpp7L13(40), cin=>outpp8L13(40), S=>outpp6L9(40) ,cout=>outpp2L9(41));
FA119L13: FA port map(A=>outpp9L13(40), B=>outpp10L13(40), cin=>outpp11L13(40), S=>outpp7L9(40) ,cout=>outpp3L9(41));
outpp8L9(40)<=outpp12L13(40);
FA120L13: FA port map(A=>outpp0L13(41), B=>outpp1L13(41), cin=>outpp2L13(41), S=>outpp4L9(41) ,cout=>outpp0L9(42));
FA121L13: FA port map(A=>outpp3L13(41), B=>outpp4L13(41), cin=>outpp5L13(41), S=>outpp5L9(41) ,cout=>outpp1L9(42));
FA122L13: FA port map(A=>outpp6L13(41), B=>outpp7L13(41), cin=>outpp8L13(41), S=>outpp6L9(41) ,cout=>outpp2L9(42));
FA123L13: FA port map(A=>outpp9L13(41), B=>outpp10L13(41), cin=>outpp11L13(41), S=>outpp7L9(41) ,cout=>outpp3L9(42));
outpp8L9(41)<=outpp12L13(41);
FA124L13: FA port map(A=>outpp0L13(42), B=>outpp1L13(42), cin=>outpp2L13(42), S=>outpp4L9(42) ,cout=>outpp0L9(43));
FA125L13: FA port map(A=>outpp3L13(42), B=>outpp4L13(42), cin=>outpp5L13(42), S=>outpp5L9(42) ,cout=>outpp1L9(43));
FA126L13: FA port map(A=>outpp6L13(42), B=>outpp7L13(42), cin=>outpp8L13(42), S=>outpp6L9(42) ,cout=>outpp2L9(43));
FA127L13: FA port map(A=>outpp9L13(42), B=>outpp10L13(42), cin=>outpp11L13(42), S=>outpp7L9(42) ,cout=>outpp3L9(43));
outpp8L9(42)<=outpp12L13(42);
FA128L13: FA port map(A=>outpp0L13(43), B=>outpp1L13(43), cin=>outpp2L13(43), S=>outpp4L9(43) ,cout=>outpp0L9(44));
FA129L13: FA port map(A=>outpp3L13(43), B=>outpp4L13(43), cin=>outpp5L13(43), S=>outpp5L9(43) ,cout=>outpp1L9(44));
FA130L13: FA port map(A=>outpp6L13(43), B=>outpp7L13(43), cin=>outpp8L13(43), S=>outpp6L9(43) ,cout=>outpp2L9(44));
FA131L13: FA port map(A=>outpp9L13(43), B=>outpp10L13(43), cin=>outpp11L13(43), S=>outpp7L9(43) ,cout=>outpp3L9(44));
outpp8L9(43)<=outpp12L13(43);
HA20L13: HA port map( A=>outpp0L13(44), B=>outpp1L13(44), S=>outpp4L9(44) ,cout=>outpp0L9(45));
FA132L13: FA port map(A=>outpp2L13(44), B=>outpp3L13(44), cin=>outpp4L13(44), S=>outpp5L9(44) ,cout=>outpp1L9(45));
FA133L13: FA port map(A=>outpp5L13(44), B=>outpp6L13(44), cin=>outpp7L13(44), S=>outpp6L9(44) ,cout=>outpp2L9(45));
FA134L13: FA port map(A=>outpp8L13(44), B=>outpp9L13(44), cin=>outpp10L13(44), S=>outpp7L9(44) ,cout=>outpp3L9(45));
outpp8L9(44)<=outpp11L13(44);
FA135L13: FA port map(A=>outpp0L13(45), B=>outpp1L13(45), cin=>outpp2L13(45), S=>outpp4L9(45) ,cout=>outpp0L9(46));
FA136L13: FA port map(A=>outpp3L13(45), B=>outpp4L13(45), cin=>outpp5L13(45), S=>outpp5L9(45) ,cout=>outpp1L9(46));
FA137L13: FA port map(A=>outpp6L13(45), B=>outpp7L13(45), cin=>outpp8L13(45), S=>outpp6L9(45) ,cout=>outpp2L9(46));
outpp7L9(45)<=outpp9L13(45);
outpp8L9(45)<=outpp10L13(45);
HA21L13: HA port map( A=>outpp0L13(46), B=>outpp1L13(46), S=>outpp3L9(46) ,cout=>outpp0L9(47));
FA138L13: FA port map(A=>outpp2L13(46), B=>outpp3L13(46), cin=>outpp4L13(46), S=>outpp4L9(46) ,cout=>outpp1L9(47));
FA139L13: FA port map(A=>outpp5L13(46), B=>outpp6L13(46), cin=>outpp7L13(46), S=>outpp5L9(46) ,cout=>outpp2L9(47));
outpp6L9(46)<=outpp8L13(46);
outpp7L9(46)<=outpp9L13(46);
outpp8L9(46)<=outpp10L13(46);
FA140L13: FA port map(A=>outpp0L13(47), B=>outpp1L13(47), cin=>outpp2L13(47), S=>outpp3L9(47) ,cout=>outpp0L9(48));
FA141L13: FA port map(A=>outpp3L13(47), B=>outpp4L13(47), cin=>outpp5L13(47), S=>outpp4L9(47) ,cout=>outpp1L9(48));
outpp5L9(47)<=outpp6L13(47);
outpp6L9(47)<=outpp7L13(47);
outpp7L9(47)<=outpp8L13(47);
outpp8L9(47)<=outpp9L13(47);
HA22L13: HA port map( A=>outpp0L13(48), B=>outpp1L13(48), S=>outpp2L9(48) ,cout=>outpp0L9(49));
FA142L13: FA port map(A=>outpp2L13(48), B=>outpp3L13(48), cin=>outpp4L13(48), S=>outpp3L9(48) ,cout=>outpp1L9(49));
outpp4L9(48)<=outpp5L13(48);
outpp5L9(48)<=outpp6L13(48);
outpp6L9(48)<=outpp7L13(48);
outpp7L9(48)<=outpp8L13(48);
outpp8L9(48)<=outpp9L13(48);
FA143L13: FA port map(A=>outpp0L13(49), B=>outpp1L13(49), cin=>outpp2L13(49), S=>outpp2L9(49) ,cout=>outpp0L9(50));
outpp3L9(49)<=outpp3L13(49);
outpp4L9(49)<=outpp4L13(49);
outpp5L9(49)<=outpp5L13(49);
outpp6L9(49)<=outpp6L13(49);
outpp7L9(49)<=outpp7L13(49);
outpp8L9(49)<=outpp8L13(49);
HA23L13: HA port map( A=>outpp0L13(50), B=>outpp1L13(50), S=>outpp1L9(50) ,cout=>outpp0L9(51));
outpp2L9(50)<=outpp2L13(50);
outpp3L9(50)<=outpp3L13(50);
outpp4L9(50)<=outpp4L13(50);
outpp5L9(50)<=outpp5L13(50);
outpp6L9(50)<=outpp6L13(50);
outpp7L9(50)<=outpp7L13(50);
outpp8L9(50)<=outpp8L13(50);
outpp1L9(51)<=outpp0L13(51);
outpp2L9(51)<=outpp1L13(51);
outpp3L9(51)<=outpp2L13(51);
outpp4L9(51)<=outpp3L13(51);
outpp5L9(51)<=outpp4L13(51);
outpp6L9(51)<=outpp5L13(51);
outpp7L9(51)<=outpp6L13(51);
outpp8L9(51)<=outpp7L13(51);
outpp0L9(52)<=outpp0L13(52);
outpp1L9(52)<=outpp1L13(52);
outpp2L9(52)<=outpp2L13(52);
outpp3L9(52)<=outpp3L13(52);
outpp4L9(52)<=outpp4L13(52);
outpp5L9(52)<=outpp5L13(52);
outpp6L9(52)<=outpp6L13(52);
outpp7L9(52)<=outpp7L13(52);
outpp8L9(52)<=outpp8L13(52);
outpp0L9(53)<=outpp0L13(53);
outpp1L9(53)<=outpp1L13(53);
outpp2L9(53)<=outpp2L13(53);
outpp3L9(53)<=outpp3L13(53);
outpp4L9(53)<=outpp4L13(53);
outpp5L9(53)<=outpp5L13(53);
outpp6L9(53)<=outpp6L13(53);
outpp7L9(53)<=outpp7L13(53);
outpp8L9(53)<=outpp8L13(53);
outpp0L9(54)<=outpp0L13(54);
outpp1L9(54)<=outpp1L13(54);
outpp2L9(54)<=outpp2L13(54);
outpp3L9(54)<=outpp3L13(54);
outpp4L9(54)<=outpp4L13(54);
outpp5L9(54)<=outpp5L13(54);
outpp6L9(54)<=outpp6L13(54);
outpp7L9(54)<=outpp7L13(54);
outpp8L9(54)<=outpp8L13(54);
outpp0L9(55)<=outpp0L13(55);
outpp1L9(55)<=outpp1L13(55);
outpp2L9(55)<=outpp2L13(55);
outpp3L9(55)<=outpp3L13(55);
outpp4L9(55)<=outpp4L13(55);
outpp5L9(55)<=outpp5L13(55);
outpp6L9(55)<=outpp6L13(55);
outpp7L9(55)<=outpp7L13(55);
outpp8L9(55)<=outpp8L13(55);
outpp0L9(56)<=outpp0L13(56);
outpp1L9(56)<=outpp1L13(56);
outpp2L9(56)<=outpp2L13(56);
outpp3L9(56)<=outpp3L13(56);
outpp4L9(56)<=outpp4L13(56);
outpp5L9(56)<=outpp5L13(56);
outpp6L9(56)<=outpp6L13(56);
outpp7L9(56)<=outpp7L13(56);
outpp8L9(56)<=outpp8L13(56);
outpp0L9(57)<=outpp0L13(57);
outpp1L9(57)<=outpp1L13(57);
outpp2L9(57)<=outpp2L13(57);
outpp3L9(57)<=outpp3L13(57);
outpp4L9(57)<=outpp4L13(57);
outpp5L9(57)<=outpp5L13(57);
outpp6L9(57)<=outpp6L13(57);
outpp7L9(57)<=outpp7L13(57);
outpp8L9(57)<=outpp8L13(57);
outpp0L9(58)<=outpp0L13(58);
outpp1L9(58)<=outpp1L13(58);
outpp2L9(58)<=outpp2L13(58);
outpp3L9(58)<=outpp3L13(58);
outpp4L9(58)<=outpp4L13(58);
outpp5L9(58)<=outpp5L13(58);
outpp6L9(58)<=outpp6L13(58);
outpp7L9(58)<=outpp7L13(58);
outpp8L9(58)<=outpp8L13(58);
outpp0L9(59)<=outpp0L13(59);
outpp1L9(59)<=outpp1L13(59);
outpp2L9(59)<=outpp2L13(59);
outpp3L9(59)<=outpp3L13(59);
outpp4L9(59)<=outpp4L13(59);
outpp5L9(59)<=outpp5L13(59);
outpp6L9(59)<=outpp6L13(59);
outpp7L9(59)<=outpp7L13(59);
outpp8L9(59)<=outpp8L13(59);
outpp0L9(60)<=outpp0L13(60);
outpp1L9(60)<=outpp1L13(60);
outpp2L9(60)<=outpp2L13(60);
outpp3L9(60)<=outpp3L13(60);
outpp4L9(60)<=outpp4L13(60);
outpp5L9(60)<=outpp5L13(60);
outpp6L9(60)<=outpp6L13(60);
outpp7L9(60)<=outpp7L13(60);
outpp8L9(60)<=outpp8L13(60);
outpp0L9(61)<=outpp0L13(61);
outpp1L9(61)<=outpp1L13(61);
outpp2L9(61)<=outpp2L13(61);
outpp3L9(61)<=outpp3L13(61);
outpp4L9(61)<=outpp4L13(61);
outpp5L9(61)<=outpp5L13(61);
outpp6L9(61)<=outpp6L13(61);
outpp7L9(61)<=outpp7L13(61);
outpp8L9(61)<=outpp8L13(61);
outpp0L9(62)<=outpp0L13(62);
outpp1L9(62)<=outpp1L13(62);
outpp2L9(62)<=outpp2L13(62);
outpp3L9(62)<=outpp3L13(62);
outpp4L9(62)<=outpp4L13(62);
outpp5L9(62)<=outpp5L13(62);
outpp6L9(62)<=outpp6L13(62);
outpp7L9(62)<=outpp7L13(62);
outpp8L9(62)<=outpp8L13(62);
outpp0L9(63)<=outpp0L13(63);
outpp1L9(63)<=outpp1L13(63);
outpp2L9(63)<=outpp2L13(63);
outpp3L9(63)<=outpp3L13(63);
outpp4L9(63)<=outpp4L13(63);
outpp5L9(63)<=outpp5L13(63);
outpp6L9(63)<=outpp6L13(63);
outpp7L9(63)<=outpp7L13(63);
outpp8L9(63)<=outpp8L13(63);
outpp0L6(0)<=outpp0L9(0);
outpp1L6(0)<=outpp1L9(0);
outpp2L6(0)<=outpp2L9(0);
outpp3L6(0)<=outpp3L9(0);
outpp4L6(0)<=outpp4L9(0);
outpp5L6(0)<=outpp5L9(0);
outpp0L6(1)<=outpp0L9(1);
outpp1L6(1)<=outpp1L9(1);
outpp2L6(1)<=outpp2L9(1);
outpp3L6(1)<=outpp3L9(1);
outpp4L6(1)<=outpp4L9(1);
outpp5L6(1)<=outpp5L9(1);
outpp0L6(2)<=outpp0L9(2);
outpp1L6(2)<=outpp1L9(2);
outpp2L6(2)<=outpp2L9(2);
outpp3L6(2)<=outpp3L9(2);
outpp4L6(2)<=outpp4L9(2);
outpp5L6(2)<=outpp5L9(2);
outpp0L6(3)<=outpp0L9(3);
outpp1L6(3)<=outpp1L9(3);
outpp2L6(3)<=outpp2L9(3);
outpp3L6(3)<=outpp3L9(3);
outpp4L6(3)<=outpp4L9(3);
outpp5L6(3)<=outpp5L9(3);
outpp0L6(4)<=outpp0L9(4);
outpp1L6(4)<=outpp1L9(4);
outpp2L6(4)<=outpp2L9(4);
outpp3L6(4)<=outpp3L9(4);
outpp4L6(4)<=outpp4L9(4);
outpp5L6(4)<=outpp5L9(4);
outpp0L6(5)<=outpp0L9(5);
outpp1L6(5)<=outpp1L9(5);
outpp2L6(5)<=outpp2L9(5);
outpp3L6(5)<=outpp3L9(5);
outpp4L6(5)<=outpp4L9(5);
outpp5L6(5)<=outpp5L9(5);
outpp0L6(6)<=outpp0L9(6);
outpp1L6(6)<=outpp1L9(6);
outpp2L6(6)<=outpp2L9(6);
outpp3L6(6)<=outpp3L9(6);
outpp4L6(6)<=outpp4L9(6);
outpp5L6(6)<=outpp5L9(6);
outpp0L6(7)<=outpp0L9(7);
outpp1L6(7)<=outpp1L9(7);
outpp2L6(7)<=outpp2L9(7);
outpp3L6(7)<=outpp3L9(7);
outpp4L6(7)<=outpp4L9(7);
outpp5L6(7)<=outpp5L9(7);
outpp0L6(8)<=outpp0L9(8);
outpp1L6(8)<=outpp1L9(8);
outpp2L6(8)<=outpp2L9(8);
outpp3L6(8)<=outpp3L9(8);
outpp4L6(8)<=outpp4L9(8);
outpp5L6(8)<=outpp5L9(8);
outpp0L6(9)<=outpp0L9(9);
outpp1L6(9)<=outpp1L9(9);
outpp2L6(9)<=outpp2L9(9);
outpp3L6(9)<=outpp3L9(9);
outpp4L6(9)<=outpp4L9(9);
outpp5L6(9)<=outpp5L9(9);
HA24L9: HA port map( A=>outpp0L9(10), B=>outpp1L9(10), S=>outpp0L6(10) ,cout=>outpp0L6(11));
outpp1L6(10)<=outpp2L9(10);
outpp2L6(10)<=outpp3L9(10);
outpp3L6(10)<=outpp4L9(10);
outpp4L6(10)<=outpp5L9(10);
outpp5L6(10)<=outpp6L9(10);
HA25L9: HA port map( A=>outpp0L9(11), B=>outpp1L9(11), S=>outpp1L6(11) ,cout=>outpp0L6(12));
outpp2L6(11)<=outpp2L9(11);
outpp3L6(11)<=outpp3L9(11);
outpp4L6(11)<=outpp4L9(11);
outpp5L6(11)<=outpp5L9(11);
HA26L9: HA port map( A=>outpp0L9(12), B=>outpp1L9(12), S=>outpp1L6(12) ,cout=>outpp0L6(13));
FA144L9: FA port map(A=>outpp2L9(12), B=>outpp3L9(12), cin=>outpp4L9(12), S=>outpp2L6(12) ,cout=>outpp1L6(13));
outpp3L6(12)<=outpp5L9(12);
outpp4L6(12)<=outpp6L9(12);
outpp5L6(12)<=outpp7L9(12);
HA27L9: HA port map( A=>outpp0L9(13), B=>outpp1L9(13), S=>outpp2L6(13) ,cout=>outpp0L6(14));
FA145L9: FA port map(A=>outpp2L9(13), B=>outpp3L9(13), cin=>outpp4L9(13), S=>outpp3L6(13) ,cout=>outpp1L6(14));
outpp4L6(13)<=outpp5L9(13);
outpp5L6(13)<=outpp6L9(13);
HA28L9: HA port map( A=>outpp0L9(14), B=>outpp1L9(14), S=>outpp2L6(14) ,cout=>outpp0L6(15));
FA146L9: FA port map(A=>outpp2L9(14), B=>outpp3L9(14), cin=>outpp4L9(14), S=>outpp3L6(14) ,cout=>outpp1L6(15));
FA147L9: FA port map(A=>outpp5L9(14), B=>outpp6L9(14), cin=>outpp7L9(14), S=>outpp4L6(14) ,cout=>outpp2L6(15));
outpp5L6(14)<=outpp8L9(14);
HA29L9: HA port map( A=>outpp0L9(15), B=>outpp1L9(15), S=>outpp3L6(15) ,cout=>outpp0L6(16));
FA148L9: FA port map(A=>outpp2L9(15), B=>outpp3L9(15), cin=>outpp4L9(15), S=>outpp4L6(15) ,cout=>outpp1L6(16));
FA149L9: FA port map(A=>outpp5L9(15), B=>outpp6L9(15), cin=>outpp7L9(15), S=>outpp5L6(15) ,cout=>outpp2L6(16));
FA150L9: FA port map(A=>outpp0L9(16), B=>outpp1L9(16), cin=>outpp2L9(16), S=>outpp3L6(16) ,cout=>outpp0L6(17));
FA151L9: FA port map(A=>outpp3L9(16), B=>outpp4L9(16), cin=>outpp5L9(16), S=>outpp4L6(16) ,cout=>outpp1L6(17));
FA152L9: FA port map(A=>outpp6L9(16), B=>outpp7L9(16), cin=>outpp8L9(16), S=>outpp5L6(16) ,cout=>outpp2L6(17));
FA153L9: FA port map(A=>outpp0L9(17), B=>outpp1L9(17), cin=>outpp2L9(17), S=>outpp3L6(17) ,cout=>outpp0L6(18));
FA154L9: FA port map(A=>outpp3L9(17), B=>outpp4L9(17), cin=>outpp5L9(17), S=>outpp4L6(17) ,cout=>outpp1L6(18));
FA155L9: FA port map(A=>outpp6L9(17), B=>outpp7L9(17), cin=>outpp8L9(17), S=>outpp5L6(17) ,cout=>outpp2L6(18));
FA156L9: FA port map(A=>outpp0L9(18), B=>outpp1L9(18), cin=>outpp2L9(18), S=>outpp3L6(18) ,cout=>outpp0L6(19));
FA157L9: FA port map(A=>outpp3L9(18), B=>outpp4L9(18), cin=>outpp5L9(18), S=>outpp4L6(18) ,cout=>outpp1L6(19));
FA158L9: FA port map(A=>outpp6L9(18), B=>outpp7L9(18), cin=>outpp8L9(18), S=>outpp5L6(18) ,cout=>outpp2L6(19));
FA159L9: FA port map(A=>outpp0L9(19), B=>outpp1L9(19), cin=>outpp2L9(19), S=>outpp3L6(19) ,cout=>outpp0L6(20));
FA160L9: FA port map(A=>outpp3L9(19), B=>outpp4L9(19), cin=>outpp5L9(19), S=>outpp4L6(19) ,cout=>outpp1L6(20));
FA161L9: FA port map(A=>outpp6L9(19), B=>outpp7L9(19), cin=>outpp8L9(19), S=>outpp5L6(19) ,cout=>outpp2L6(20));
FA162L9: FA port map(A=>outpp0L9(20), B=>outpp1L9(20), cin=>outpp2L9(20), S=>outpp3L6(20) ,cout=>outpp0L6(21));
FA163L9: FA port map(A=>outpp3L9(20), B=>outpp4L9(20), cin=>outpp5L9(20), S=>outpp4L6(20) ,cout=>outpp1L6(21));
FA164L9: FA port map(A=>outpp6L9(20), B=>outpp7L9(20), cin=>outpp8L9(20), S=>outpp5L6(20) ,cout=>outpp2L6(21));
FA165L9: FA port map(A=>outpp0L9(21), B=>outpp1L9(21), cin=>outpp2L9(21), S=>outpp3L6(21) ,cout=>outpp0L6(22));
FA166L9: FA port map(A=>outpp3L9(21), B=>outpp4L9(21), cin=>outpp5L9(21), S=>outpp4L6(21) ,cout=>outpp1L6(22));
FA167L9: FA port map(A=>outpp6L9(21), B=>outpp7L9(21), cin=>outpp8L9(21), S=>outpp5L6(21) ,cout=>outpp2L6(22));
FA168L9: FA port map(A=>outpp0L9(22), B=>outpp1L9(22), cin=>outpp2L9(22), S=>outpp3L6(22) ,cout=>outpp0L6(23));
FA169L9: FA port map(A=>outpp3L9(22), B=>outpp4L9(22), cin=>outpp5L9(22), S=>outpp4L6(22) ,cout=>outpp1L6(23));
FA170L9: FA port map(A=>outpp6L9(22), B=>outpp7L9(22), cin=>outpp8L9(22), S=>outpp5L6(22) ,cout=>outpp2L6(23));
FA171L9: FA port map(A=>outpp0L9(23), B=>outpp1L9(23), cin=>outpp2L9(23), S=>outpp3L6(23) ,cout=>outpp0L6(24));
FA172L9: FA port map(A=>outpp3L9(23), B=>outpp4L9(23), cin=>outpp5L9(23), S=>outpp4L6(23) ,cout=>outpp1L6(24));
FA173L9: FA port map(A=>outpp6L9(23), B=>outpp7L9(23), cin=>outpp8L9(23), S=>outpp5L6(23) ,cout=>outpp2L6(24));
FA174L9: FA port map(A=>outpp0L9(24), B=>outpp1L9(24), cin=>outpp2L9(24), S=>outpp3L6(24) ,cout=>outpp0L6(25));
FA175L9: FA port map(A=>outpp3L9(24), B=>outpp4L9(24), cin=>outpp5L9(24), S=>outpp4L6(24) ,cout=>outpp1L6(25));
FA176L9: FA port map(A=>outpp6L9(24), B=>outpp7L9(24), cin=>outpp8L9(24), S=>outpp5L6(24) ,cout=>outpp2L6(25));
FA177L9: FA port map(A=>outpp0L9(25), B=>outpp1L9(25), cin=>outpp2L9(25), S=>outpp3L6(25) ,cout=>outpp0L6(26));
FA178L9: FA port map(A=>outpp3L9(25), B=>outpp4L9(25), cin=>outpp5L9(25), S=>outpp4L6(25) ,cout=>outpp1L6(26));
FA179L9: FA port map(A=>outpp6L9(25), B=>outpp7L9(25), cin=>outpp8L9(25), S=>outpp5L6(25) ,cout=>outpp2L6(26));
FA180L9: FA port map(A=>outpp0L9(26), B=>outpp1L9(26), cin=>outpp2L9(26), S=>outpp3L6(26) ,cout=>outpp0L6(27));
FA181L9: FA port map(A=>outpp3L9(26), B=>outpp4L9(26), cin=>outpp5L9(26), S=>outpp4L6(26) ,cout=>outpp1L6(27));
FA182L9: FA port map(A=>outpp6L9(26), B=>outpp7L9(26), cin=>outpp8L9(26), S=>outpp5L6(26) ,cout=>outpp2L6(27));
FA183L9: FA port map(A=>outpp0L9(27), B=>outpp1L9(27), cin=>outpp2L9(27), S=>outpp3L6(27) ,cout=>outpp0L6(28));
FA184L9: FA port map(A=>outpp3L9(27), B=>outpp4L9(27), cin=>outpp5L9(27), S=>outpp4L6(27) ,cout=>outpp1L6(28));
FA185L9: FA port map(A=>outpp6L9(27), B=>outpp7L9(27), cin=>outpp8L9(27), S=>outpp5L6(27) ,cout=>outpp2L6(28));
FA186L9: FA port map(A=>outpp0L9(28), B=>outpp1L9(28), cin=>outpp2L9(28), S=>outpp3L6(28) ,cout=>outpp0L6(29));
FA187L9: FA port map(A=>outpp3L9(28), B=>outpp4L9(28), cin=>outpp5L9(28), S=>outpp4L6(28) ,cout=>outpp1L6(29));
FA188L9: FA port map(A=>outpp6L9(28), B=>outpp7L9(28), cin=>outpp8L9(28), S=>outpp5L6(28) ,cout=>outpp2L6(29));
FA189L9: FA port map(A=>outpp0L9(29), B=>outpp1L9(29), cin=>outpp2L9(29), S=>outpp3L6(29) ,cout=>outpp0L6(30));
FA190L9: FA port map(A=>outpp3L9(29), B=>outpp4L9(29), cin=>outpp5L9(29), S=>outpp4L6(29) ,cout=>outpp1L6(30));
FA191L9: FA port map(A=>outpp6L9(29), B=>outpp7L9(29), cin=>outpp8L9(29), S=>outpp5L6(29) ,cout=>outpp2L6(30));
FA192L9: FA port map(A=>outpp0L9(30), B=>outpp1L9(30), cin=>outpp2L9(30), S=>outpp3L6(30) ,cout=>outpp0L6(31));
FA193L9: FA port map(A=>outpp3L9(30), B=>outpp4L9(30), cin=>outpp5L9(30), S=>outpp4L6(30) ,cout=>outpp1L6(31));
FA194L9: FA port map(A=>outpp6L9(30), B=>outpp7L9(30), cin=>outpp8L9(30), S=>outpp5L6(30) ,cout=>outpp2L6(31));
FA195L9: FA port map(A=>outpp0L9(31), B=>outpp1L9(31), cin=>outpp2L9(31), S=>outpp3L6(31) ,cout=>outpp0L6(32));
FA196L9: FA port map(A=>outpp3L9(31), B=>outpp4L9(31), cin=>outpp5L9(31), S=>outpp4L6(31) ,cout=>outpp1L6(32));
FA197L9: FA port map(A=>outpp6L9(31), B=>outpp7L9(31), cin=>outpp8L9(31), S=>outpp5L6(31) ,cout=>outpp2L6(32));
FA198L9: FA port map(A=>outpp0L9(32), B=>outpp1L9(32), cin=>outpp2L9(32), S=>outpp3L6(32) ,cout=>outpp0L6(33));
FA199L9: FA port map(A=>outpp3L9(32), B=>outpp4L9(32), cin=>outpp5L9(32), S=>outpp4L6(32) ,cout=>outpp1L6(33));
FA200L9: FA port map(A=>outpp6L9(32), B=>outpp7L9(32), cin=>outpp8L9(32), S=>outpp5L6(32) ,cout=>outpp2L6(33));
FA201L9: FA port map(A=>outpp0L9(33), B=>outpp1L9(33), cin=>outpp2L9(33), S=>outpp3L6(33) ,cout=>outpp0L6(34));
FA202L9: FA port map(A=>outpp3L9(33), B=>outpp4L9(33), cin=>outpp5L9(33), S=>outpp4L6(33) ,cout=>outpp1L6(34));
FA203L9: FA port map(A=>outpp6L9(33), B=>outpp7L9(33), cin=>outpp8L9(33), S=>outpp5L6(33) ,cout=>outpp2L6(34));
FA204L9: FA port map(A=>outpp0L9(34), B=>outpp1L9(34), cin=>outpp2L9(34), S=>outpp3L6(34) ,cout=>outpp0L6(35));
FA205L9: FA port map(A=>outpp3L9(34), B=>outpp4L9(34), cin=>outpp5L9(34), S=>outpp4L6(34) ,cout=>outpp1L6(35));
FA206L9: FA port map(A=>outpp6L9(34), B=>outpp7L9(34), cin=>outpp8L9(34), S=>outpp5L6(34) ,cout=>outpp2L6(35));
FA207L9: FA port map(A=>outpp0L9(35), B=>outpp1L9(35), cin=>outpp2L9(35), S=>outpp3L6(35) ,cout=>outpp0L6(36));
FA208L9: FA port map(A=>outpp3L9(35), B=>outpp4L9(35), cin=>outpp5L9(35), S=>outpp4L6(35) ,cout=>outpp1L6(36));
FA209L9: FA port map(A=>outpp6L9(35), B=>outpp7L9(35), cin=>outpp8L9(35), S=>outpp5L6(35) ,cout=>outpp2L6(36));
FA210L9: FA port map(A=>outpp0L9(36), B=>outpp1L9(36), cin=>outpp2L9(36), S=>outpp3L6(36) ,cout=>outpp0L6(37));
FA211L9: FA port map(A=>outpp3L9(36), B=>outpp4L9(36), cin=>outpp5L9(36), S=>outpp4L6(36) ,cout=>outpp1L6(37));
FA212L9: FA port map(A=>outpp6L9(36), B=>outpp7L9(36), cin=>outpp8L9(36), S=>outpp5L6(36) ,cout=>outpp2L6(37));
FA213L9: FA port map(A=>outpp0L9(37), B=>outpp1L9(37), cin=>outpp2L9(37), S=>outpp3L6(37) ,cout=>outpp0L6(38));
FA214L9: FA port map(A=>outpp3L9(37), B=>outpp4L9(37), cin=>outpp5L9(37), S=>outpp4L6(37) ,cout=>outpp1L6(38));
FA215L9: FA port map(A=>outpp6L9(37), B=>outpp7L9(37), cin=>outpp8L9(37), S=>outpp5L6(37) ,cout=>outpp2L6(38));
FA216L9: FA port map(A=>outpp0L9(38), B=>outpp1L9(38), cin=>outpp2L9(38), S=>outpp3L6(38) ,cout=>outpp0L6(39));
FA217L9: FA port map(A=>outpp3L9(38), B=>outpp4L9(38), cin=>outpp5L9(38), S=>outpp4L6(38) ,cout=>outpp1L6(39));
FA218L9: FA port map(A=>outpp6L9(38), B=>outpp7L9(38), cin=>outpp8L9(38), S=>outpp5L6(38) ,cout=>outpp2L6(39));
FA219L9: FA port map(A=>outpp0L9(39), B=>outpp1L9(39), cin=>outpp2L9(39), S=>outpp3L6(39) ,cout=>outpp0L6(40));
FA220L9: FA port map(A=>outpp3L9(39), B=>outpp4L9(39), cin=>outpp5L9(39), S=>outpp4L6(39) ,cout=>outpp1L6(40));
FA221L9: FA port map(A=>outpp6L9(39), B=>outpp7L9(39), cin=>outpp8L9(39), S=>outpp5L6(39) ,cout=>outpp2L6(40));
FA222L9: FA port map(A=>outpp0L9(40), B=>outpp1L9(40), cin=>outpp2L9(40), S=>outpp3L6(40) ,cout=>outpp0L6(41));
FA223L9: FA port map(A=>outpp3L9(40), B=>outpp4L9(40), cin=>outpp5L9(40), S=>outpp4L6(40) ,cout=>outpp1L6(41));
FA224L9: FA port map(A=>outpp6L9(40), B=>outpp7L9(40), cin=>outpp8L9(40), S=>outpp5L6(40) ,cout=>outpp2L6(41));
FA225L9: FA port map(A=>outpp0L9(41), B=>outpp1L9(41), cin=>outpp2L9(41), S=>outpp3L6(41) ,cout=>outpp0L6(42));
FA226L9: FA port map(A=>outpp3L9(41), B=>outpp4L9(41), cin=>outpp5L9(41), S=>outpp4L6(41) ,cout=>outpp1L6(42));
FA227L9: FA port map(A=>outpp6L9(41), B=>outpp7L9(41), cin=>outpp8L9(41), S=>outpp5L6(41) ,cout=>outpp2L6(42));
FA228L9: FA port map(A=>outpp0L9(42), B=>outpp1L9(42), cin=>outpp2L9(42), S=>outpp3L6(42) ,cout=>outpp0L6(43));
FA229L9: FA port map(A=>outpp3L9(42), B=>outpp4L9(42), cin=>outpp5L9(42), S=>outpp4L6(42) ,cout=>outpp1L6(43));
FA230L9: FA port map(A=>outpp6L9(42), B=>outpp7L9(42), cin=>outpp8L9(42), S=>outpp5L6(42) ,cout=>outpp2L6(43));
FA231L9: FA port map(A=>outpp0L9(43), B=>outpp1L9(43), cin=>outpp2L9(43), S=>outpp3L6(43) ,cout=>outpp0L6(44));
FA232L9: FA port map(A=>outpp3L9(43), B=>outpp4L9(43), cin=>outpp5L9(43), S=>outpp4L6(43) ,cout=>outpp1L6(44));
FA233L9: FA port map(A=>outpp6L9(43), B=>outpp7L9(43), cin=>outpp8L9(43), S=>outpp5L6(43) ,cout=>outpp2L6(44));
FA234L9: FA port map(A=>outpp0L9(44), B=>outpp1L9(44), cin=>outpp2L9(44), S=>outpp3L6(44) ,cout=>outpp0L6(45));
FA235L9: FA port map(A=>outpp3L9(44), B=>outpp4L9(44), cin=>outpp5L9(44), S=>outpp4L6(44) ,cout=>outpp1L6(45));
FA236L9: FA port map(A=>outpp6L9(44), B=>outpp7L9(44), cin=>outpp8L9(44), S=>outpp5L6(44) ,cout=>outpp2L6(45));
FA237L9: FA port map(A=>outpp0L9(45), B=>outpp1L9(45), cin=>outpp2L9(45), S=>outpp3L6(45) ,cout=>outpp0L6(46));
FA238L9: FA port map(A=>outpp3L9(45), B=>outpp4L9(45), cin=>outpp5L9(45), S=>outpp4L6(45) ,cout=>outpp1L6(46));
FA239L9: FA port map(A=>outpp6L9(45), B=>outpp7L9(45), cin=>outpp8L9(45), S=>outpp5L6(45) ,cout=>outpp2L6(46));
FA240L9: FA port map(A=>outpp0L9(46), B=>outpp1L9(46), cin=>outpp2L9(46), S=>outpp3L6(46) ,cout=>outpp0L6(47));
FA241L9: FA port map(A=>outpp3L9(46), B=>outpp4L9(46), cin=>outpp5L9(46), S=>outpp4L6(46) ,cout=>outpp1L6(47));
FA242L9: FA port map(A=>outpp6L9(46), B=>outpp7L9(46), cin=>outpp8L9(46), S=>outpp5L6(46) ,cout=>outpp2L6(47));
FA243L9: FA port map(A=>outpp0L9(47), B=>outpp1L9(47), cin=>outpp2L9(47), S=>outpp3L6(47) ,cout=>outpp0L6(48));
FA244L9: FA port map(A=>outpp3L9(47), B=>outpp4L9(47), cin=>outpp5L9(47), S=>outpp4L6(47) ,cout=>outpp1L6(48));
FA245L9: FA port map(A=>outpp6L9(47), B=>outpp7L9(47), cin=>outpp8L9(47), S=>outpp5L6(47) ,cout=>outpp2L6(48));
FA246L9: FA port map(A=>outpp0L9(48), B=>outpp1L9(48), cin=>outpp2L9(48), S=>outpp3L6(48) ,cout=>outpp0L6(49));
FA247L9: FA port map(A=>outpp3L9(48), B=>outpp4L9(48), cin=>outpp5L9(48), S=>outpp4L6(48) ,cout=>outpp1L6(49));
FA248L9: FA port map(A=>outpp6L9(48), B=>outpp7L9(48), cin=>outpp8L9(48), S=>outpp5L6(48) ,cout=>outpp2L6(49));
FA249L9: FA port map(A=>outpp0L9(49), B=>outpp1L9(49), cin=>outpp2L9(49), S=>outpp3L6(49) ,cout=>outpp0L6(50));
FA250L9: FA port map(A=>outpp3L9(49), B=>outpp4L9(49), cin=>outpp5L9(49), S=>outpp4L6(49) ,cout=>outpp1L6(50));
FA251L9: FA port map(A=>outpp6L9(49), B=>outpp7L9(49), cin=>outpp8L9(49), S=>outpp5L6(49) ,cout=>outpp2L6(50));
FA252L9: FA port map(A=>outpp0L9(50), B=>outpp1L9(50), cin=>outpp2L9(50), S=>outpp3L6(50) ,cout=>outpp0L6(51));
FA253L9: FA port map(A=>outpp3L9(50), B=>outpp4L9(50), cin=>outpp5L9(50), S=>outpp4L6(50) ,cout=>outpp1L6(51));
FA254L9: FA port map(A=>outpp6L9(50), B=>outpp7L9(50), cin=>outpp8L9(50), S=>outpp5L6(50) ,cout=>outpp2L6(51));
FA255L9: FA port map(A=>outpp0L9(51), B=>outpp1L9(51), cin=>outpp2L9(51), S=>outpp3L6(51) ,cout=>outpp0L6(52));
FA256L9: FA port map(A=>outpp3L9(51), B=>outpp4L9(51), cin=>outpp5L9(51), S=>outpp4L6(51) ,cout=>outpp1L6(52));
FA257L9: FA port map(A=>outpp6L9(51), B=>outpp7L9(51), cin=>outpp8L9(51), S=>outpp5L6(51) ,cout=>outpp2L6(52));
HA30L9: HA port map( A=>outpp0L9(52), B=>outpp1L9(52), S=>outpp3L6(52) ,cout=>outpp0L6(53));
FA258L9: FA port map(A=>outpp2L9(52), B=>outpp3L9(52), cin=>outpp4L9(52), S=>outpp4L6(52) ,cout=>outpp1L6(53));
FA259L9: FA port map(A=>outpp5L9(52), B=>outpp6L9(52), cin=>outpp7L9(52), S=>outpp5L6(52) ,cout=>outpp2L6(53));
FA260L9: FA port map(A=>outpp0L9(53), B=>outpp1L9(53), cin=>outpp2L9(53), S=>outpp3L6(53) ,cout=>outpp0L6(54));
FA261L9: FA port map(A=>outpp3L9(53), B=>outpp4L9(53), cin=>outpp5L9(53), S=>outpp4L6(53) ,cout=>outpp1L6(54));
outpp5L6(53)<=outpp6L9(53);
HA31L9: HA port map( A=>outpp0L9(54), B=>outpp1L9(54), S=>outpp2L6(54) ,cout=>outpp0L6(55));
FA262L9: FA port map(A=>outpp2L9(54), B=>outpp3L9(54), cin=>outpp4L9(54), S=>outpp3L6(54) ,cout=>outpp1L6(55));
outpp4L6(54)<=outpp5L9(54);
outpp5L6(54)<=outpp6L9(54);
FA263L9: FA port map(A=>outpp0L9(55), B=>outpp1L9(55), cin=>outpp2L9(55), S=>outpp2L6(55) ,cout=>outpp0L6(56));
outpp3L6(55)<=outpp3L9(55);
outpp4L6(55)<=outpp4L9(55);
outpp5L6(55)<=outpp5L9(55);
HA32L9: HA port map( A=>outpp0L9(56), B=>outpp1L9(56), S=>outpp1L6(56) ,cout=>outpp0L6(57));
outpp2L6(56)<=outpp2L9(56);
outpp3L6(56)<=outpp3L9(56);
outpp4L6(56)<=outpp4L9(56);
outpp5L6(56)<=outpp5L9(56);
outpp1L6(57)<=outpp0L9(57);
outpp2L6(57)<=outpp1L9(57);
outpp3L6(57)<=outpp2L9(57);
outpp4L6(57)<=outpp3L9(57);
outpp5L6(57)<=outpp4L9(57);
outpp0L6(58)<=outpp0L9(58);
outpp1L6(58)<=outpp1L9(58);
outpp2L6(58)<=outpp2L9(58);
outpp3L6(58)<=outpp3L9(58);
outpp4L6(58)<=outpp4L9(58);
outpp5L6(58)<=outpp5L9(58);
outpp0L6(59)<=outpp0L9(59);
outpp1L6(59)<=outpp1L9(59);
outpp2L6(59)<=outpp2L9(59);
outpp3L6(59)<=outpp3L9(59);
outpp4L6(59)<=outpp4L9(59);
outpp5L6(59)<=outpp5L9(59);
outpp0L6(60)<=outpp0L9(60);
outpp1L6(60)<=outpp1L9(60);
outpp2L6(60)<=outpp2L9(60);
outpp3L6(60)<=outpp3L9(60);
outpp4L6(60)<=outpp4L9(60);
outpp5L6(60)<=outpp5L9(60);
outpp0L6(61)<=outpp0L9(61);
outpp1L6(61)<=outpp1L9(61);
outpp2L6(61)<=outpp2L9(61);
outpp3L6(61)<=outpp3L9(61);
outpp4L6(61)<=outpp4L9(61);
outpp5L6(61)<=outpp5L9(61);
outpp0L6(62)<=outpp0L9(62);
outpp1L6(62)<=outpp1L9(62);
outpp2L6(62)<=outpp2L9(62);
outpp3L6(62)<=outpp3L9(62);
outpp4L6(62)<=outpp4L9(62);
outpp5L6(62)<=outpp5L9(62);
outpp0L6(63)<=outpp0L9(63);
outpp1L6(63)<=outpp1L9(63);
outpp2L6(63)<=outpp2L9(63);
outpp3L6(63)<=outpp3L9(63);
outpp4L6(63)<=outpp4L9(63);
outpp5L6(63)<=outpp5L9(63);
outpp0L4(0)<=outpp0L6(0);
outpp1L4(0)<=outpp1L6(0);
outpp2L4(0)<=outpp2L6(0);
outpp3L4(0)<=outpp3L6(0);
outpp0L4(1)<=outpp0L6(1);
outpp1L4(1)<=outpp1L6(1);
outpp2L4(1)<=outpp2L6(1);
outpp3L4(1)<=outpp3L6(1);
outpp0L4(2)<=outpp0L6(2);
outpp1L4(2)<=outpp1L6(2);
outpp2L4(2)<=outpp2L6(2);
outpp3L4(2)<=outpp3L6(2);
outpp0L4(3)<=outpp0L6(3);
outpp1L4(3)<=outpp1L6(3);
outpp2L4(3)<=outpp2L6(3);
outpp3L4(3)<=outpp3L6(3);
outpp0L4(4)<=outpp0L6(4);
outpp1L4(4)<=outpp1L6(4);
outpp2L4(4)<=outpp2L6(4);
outpp3L4(4)<=outpp3L6(4);
outpp0L4(5)<=outpp0L6(5);
outpp1L4(5)<=outpp1L6(5);
outpp2L4(5)<=outpp2L6(5);
outpp3L4(5)<=outpp3L6(5);
HA33L6: HA port map( A=>outpp0L6(6), B=>outpp1L6(6), S=>outpp0L4(6) ,cout=>outpp0L4(7));
outpp1L4(6)<=outpp2L6(6);
outpp2L4(6)<=outpp3L6(6);
outpp3L4(6)<=outpp4L6(6);
HA34L6: HA port map( A=>outpp0L6(7), B=>outpp1L6(7), S=>outpp1L4(7) ,cout=>outpp0L4(8));
outpp2L4(7)<=outpp2L6(7);
outpp3L4(7)<=outpp3L6(7);
HA35L6: HA port map( A=>outpp0L6(8), B=>outpp1L6(8), S=>outpp1L4(8) ,cout=>outpp0L4(9));
FA264L6: FA port map(A=>outpp2L6(8), B=>outpp3L6(8), cin=>outpp4L6(8), S=>outpp2L4(8) ,cout=>outpp1L4(9));
outpp3L4(8)<=outpp5L6(8);
HA36L6: HA port map( A=>outpp0L6(9), B=>outpp1L6(9), S=>outpp2L4(9) ,cout=>outpp0L4(10));
FA265L6: FA port map(A=>outpp2L6(9), B=>outpp3L6(9), cin=>outpp4L6(9), S=>outpp3L4(9) ,cout=>outpp1L4(10));
FA266L6: FA port map(A=>outpp0L6(10), B=>outpp1L6(10), cin=>outpp2L6(10), S=>outpp2L4(10) ,cout=>outpp0L4(11));
FA267L6: FA port map(A=>outpp3L6(10), B=>outpp4L6(10), cin=>outpp5L6(10), S=>outpp3L4(10) ,cout=>outpp1L4(11));
FA268L6: FA port map(A=>outpp0L6(11), B=>outpp1L6(11), cin=>outpp2L6(11), S=>outpp2L4(11) ,cout=>outpp0L4(12));
FA269L6: FA port map(A=>outpp3L6(11), B=>outpp4L6(11), cin=>outpp5L6(11), S=>outpp3L4(11) ,cout=>outpp1L4(12));
FA270L6: FA port map(A=>outpp0L6(12), B=>outpp1L6(12), cin=>outpp2L6(12), S=>outpp2L4(12) ,cout=>outpp0L4(13));
FA271L6: FA port map(A=>outpp3L6(12), B=>outpp4L6(12), cin=>outpp5L6(12), S=>outpp3L4(12) ,cout=>outpp1L4(13));
FA272L6: FA port map(A=>outpp0L6(13), B=>outpp1L6(13), cin=>outpp2L6(13), S=>outpp2L4(13) ,cout=>outpp0L4(14));
FA273L6: FA port map(A=>outpp3L6(13), B=>outpp4L6(13), cin=>outpp5L6(13), S=>outpp3L4(13) ,cout=>outpp1L4(14));
FA274L6: FA port map(A=>outpp0L6(14), B=>outpp1L6(14), cin=>outpp2L6(14), S=>outpp2L4(14) ,cout=>outpp0L4(15));
FA275L6: FA port map(A=>outpp3L6(14), B=>outpp4L6(14), cin=>outpp5L6(14), S=>outpp3L4(14) ,cout=>outpp1L4(15));
FA276L6: FA port map(A=>outpp0L6(15), B=>outpp1L6(15), cin=>outpp2L6(15), S=>outpp2L4(15) ,cout=>outpp0L4(16));
FA277L6: FA port map(A=>outpp3L6(15), B=>outpp4L6(15), cin=>outpp5L6(15), S=>outpp3L4(15) ,cout=>outpp1L4(16));
FA278L6: FA port map(A=>outpp0L6(16), B=>outpp1L6(16), cin=>outpp2L6(16), S=>outpp2L4(16) ,cout=>outpp0L4(17));
FA279L6: FA port map(A=>outpp3L6(16), B=>outpp4L6(16), cin=>outpp5L6(16), S=>outpp3L4(16) ,cout=>outpp1L4(17));
FA280L6: FA port map(A=>outpp0L6(17), B=>outpp1L6(17), cin=>outpp2L6(17), S=>outpp2L4(17) ,cout=>outpp0L4(18));
FA281L6: FA port map(A=>outpp3L6(17), B=>outpp4L6(17), cin=>outpp5L6(17), S=>outpp3L4(17) ,cout=>outpp1L4(18));
FA282L6: FA port map(A=>outpp0L6(18), B=>outpp1L6(18), cin=>outpp2L6(18), S=>outpp2L4(18) ,cout=>outpp0L4(19));
FA283L6: FA port map(A=>outpp3L6(18), B=>outpp4L6(18), cin=>outpp5L6(18), S=>outpp3L4(18) ,cout=>outpp1L4(19));
FA284L6: FA port map(A=>outpp0L6(19), B=>outpp1L6(19), cin=>outpp2L6(19), S=>outpp2L4(19) ,cout=>outpp0L4(20));
FA285L6: FA port map(A=>outpp3L6(19), B=>outpp4L6(19), cin=>outpp5L6(19), S=>outpp3L4(19) ,cout=>outpp1L4(20));
FA286L6: FA port map(A=>outpp0L6(20), B=>outpp1L6(20), cin=>outpp2L6(20), S=>outpp2L4(20) ,cout=>outpp0L4(21));
FA287L6: FA port map(A=>outpp3L6(20), B=>outpp4L6(20), cin=>outpp5L6(20), S=>outpp3L4(20) ,cout=>outpp1L4(21));
FA288L6: FA port map(A=>outpp0L6(21), B=>outpp1L6(21), cin=>outpp2L6(21), S=>outpp2L4(21) ,cout=>outpp0L4(22));
FA289L6: FA port map(A=>outpp3L6(21), B=>outpp4L6(21), cin=>outpp5L6(21), S=>outpp3L4(21) ,cout=>outpp1L4(22));
FA290L6: FA port map(A=>outpp0L6(22), B=>outpp1L6(22), cin=>outpp2L6(22), S=>outpp2L4(22) ,cout=>outpp0L4(23));
FA291L6: FA port map(A=>outpp3L6(22), B=>outpp4L6(22), cin=>outpp5L6(22), S=>outpp3L4(22) ,cout=>outpp1L4(23));
FA292L6: FA port map(A=>outpp0L6(23), B=>outpp1L6(23), cin=>outpp2L6(23), S=>outpp2L4(23) ,cout=>outpp0L4(24));
FA293L6: FA port map(A=>outpp3L6(23), B=>outpp4L6(23), cin=>outpp5L6(23), S=>outpp3L4(23) ,cout=>outpp1L4(24));
FA294L6: FA port map(A=>outpp0L6(24), B=>outpp1L6(24), cin=>outpp2L6(24), S=>outpp2L4(24) ,cout=>outpp0L4(25));
FA295L6: FA port map(A=>outpp3L6(24), B=>outpp4L6(24), cin=>outpp5L6(24), S=>outpp3L4(24) ,cout=>outpp1L4(25));
FA296L6: FA port map(A=>outpp0L6(25), B=>outpp1L6(25), cin=>outpp2L6(25), S=>outpp2L4(25) ,cout=>outpp0L4(26));
FA297L6: FA port map(A=>outpp3L6(25), B=>outpp4L6(25), cin=>outpp5L6(25), S=>outpp3L4(25) ,cout=>outpp1L4(26));
FA298L6: FA port map(A=>outpp0L6(26), B=>outpp1L6(26), cin=>outpp2L6(26), S=>outpp2L4(26) ,cout=>outpp0L4(27));
FA299L6: FA port map(A=>outpp3L6(26), B=>outpp4L6(26), cin=>outpp5L6(26), S=>outpp3L4(26) ,cout=>outpp1L4(27));
FA300L6: FA port map(A=>outpp0L6(27), B=>outpp1L6(27), cin=>outpp2L6(27), S=>outpp2L4(27) ,cout=>outpp0L4(28));
FA301L6: FA port map(A=>outpp3L6(27), B=>outpp4L6(27), cin=>outpp5L6(27), S=>outpp3L4(27) ,cout=>outpp1L4(28));
FA302L6: FA port map(A=>outpp0L6(28), B=>outpp1L6(28), cin=>outpp2L6(28), S=>outpp2L4(28) ,cout=>outpp0L4(29));
FA303L6: FA port map(A=>outpp3L6(28), B=>outpp4L6(28), cin=>outpp5L6(28), S=>outpp3L4(28) ,cout=>outpp1L4(29));
FA304L6: FA port map(A=>outpp0L6(29), B=>outpp1L6(29), cin=>outpp2L6(29), S=>outpp2L4(29) ,cout=>outpp0L4(30));
FA305L6: FA port map(A=>outpp3L6(29), B=>outpp4L6(29), cin=>outpp5L6(29), S=>outpp3L4(29) ,cout=>outpp1L4(30));
FA306L6: FA port map(A=>outpp0L6(30), B=>outpp1L6(30), cin=>outpp2L6(30), S=>outpp2L4(30) ,cout=>outpp0L4(31));
FA307L6: FA port map(A=>outpp3L6(30), B=>outpp4L6(30), cin=>outpp5L6(30), S=>outpp3L4(30) ,cout=>outpp1L4(31));
FA308L6: FA port map(A=>outpp0L6(31), B=>outpp1L6(31), cin=>outpp2L6(31), S=>outpp2L4(31) ,cout=>outpp0L4(32));
FA309L6: FA port map(A=>outpp3L6(31), B=>outpp4L6(31), cin=>outpp5L6(31), S=>outpp3L4(31) ,cout=>outpp1L4(32));
FA310L6: FA port map(A=>outpp0L6(32), B=>outpp1L6(32), cin=>outpp2L6(32), S=>outpp2L4(32) ,cout=>outpp0L4(33));
FA311L6: FA port map(A=>outpp3L6(32), B=>outpp4L6(32), cin=>outpp5L6(32), S=>outpp3L4(32) ,cout=>outpp1L4(33));
FA312L6: FA port map(A=>outpp0L6(33), B=>outpp1L6(33), cin=>outpp2L6(33), S=>outpp2L4(33) ,cout=>outpp0L4(34));
FA313L6: FA port map(A=>outpp3L6(33), B=>outpp4L6(33), cin=>outpp5L6(33), S=>outpp3L4(33) ,cout=>outpp1L4(34));
FA314L6: FA port map(A=>outpp0L6(34), B=>outpp1L6(34), cin=>outpp2L6(34), S=>outpp2L4(34) ,cout=>outpp0L4(35));
FA315L6: FA port map(A=>outpp3L6(34), B=>outpp4L6(34), cin=>outpp5L6(34), S=>outpp3L4(34) ,cout=>outpp1L4(35));
FA316L6: FA port map(A=>outpp0L6(35), B=>outpp1L6(35), cin=>outpp2L6(35), S=>outpp2L4(35) ,cout=>outpp0L4(36));
FA317L6: FA port map(A=>outpp3L6(35), B=>outpp4L6(35), cin=>outpp5L6(35), S=>outpp3L4(35) ,cout=>outpp1L4(36));
FA318L6: FA port map(A=>outpp0L6(36), B=>outpp1L6(36), cin=>outpp2L6(36), S=>outpp2L4(36) ,cout=>outpp0L4(37));
FA319L6: FA port map(A=>outpp3L6(36), B=>outpp4L6(36), cin=>outpp5L6(36), S=>outpp3L4(36) ,cout=>outpp1L4(37));
FA320L6: FA port map(A=>outpp0L6(37), B=>outpp1L6(37), cin=>outpp2L6(37), S=>outpp2L4(37) ,cout=>outpp0L4(38));
FA321L6: FA port map(A=>outpp3L6(37), B=>outpp4L6(37), cin=>outpp5L6(37), S=>outpp3L4(37) ,cout=>outpp1L4(38));
FA322L6: FA port map(A=>outpp0L6(38), B=>outpp1L6(38), cin=>outpp2L6(38), S=>outpp2L4(38) ,cout=>outpp0L4(39));
FA323L6: FA port map(A=>outpp3L6(38), B=>outpp4L6(38), cin=>outpp5L6(38), S=>outpp3L4(38) ,cout=>outpp1L4(39));
FA324L6: FA port map(A=>outpp0L6(39), B=>outpp1L6(39), cin=>outpp2L6(39), S=>outpp2L4(39) ,cout=>outpp0L4(40));
FA325L6: FA port map(A=>outpp3L6(39), B=>outpp4L6(39), cin=>outpp5L6(39), S=>outpp3L4(39) ,cout=>outpp1L4(40));
FA326L6: FA port map(A=>outpp0L6(40), B=>outpp1L6(40), cin=>outpp2L6(40), S=>outpp2L4(40) ,cout=>outpp0L4(41));
FA327L6: FA port map(A=>outpp3L6(40), B=>outpp4L6(40), cin=>outpp5L6(40), S=>outpp3L4(40) ,cout=>outpp1L4(41));
FA328L6: FA port map(A=>outpp0L6(41), B=>outpp1L6(41), cin=>outpp2L6(41), S=>outpp2L4(41) ,cout=>outpp0L4(42));
FA329L6: FA port map(A=>outpp3L6(41), B=>outpp4L6(41), cin=>outpp5L6(41), S=>outpp3L4(41) ,cout=>outpp1L4(42));
FA330L6: FA port map(A=>outpp0L6(42), B=>outpp1L6(42), cin=>outpp2L6(42), S=>outpp2L4(42) ,cout=>outpp0L4(43));
FA331L6: FA port map(A=>outpp3L6(42), B=>outpp4L6(42), cin=>outpp5L6(42), S=>outpp3L4(42) ,cout=>outpp1L4(43));
FA332L6: FA port map(A=>outpp0L6(43), B=>outpp1L6(43), cin=>outpp2L6(43), S=>outpp2L4(43) ,cout=>outpp0L4(44));
FA333L6: FA port map(A=>outpp3L6(43), B=>outpp4L6(43), cin=>outpp5L6(43), S=>outpp3L4(43) ,cout=>outpp1L4(44));
FA334L6: FA port map(A=>outpp0L6(44), B=>outpp1L6(44), cin=>outpp2L6(44), S=>outpp2L4(44) ,cout=>outpp0L4(45));
FA335L6: FA port map(A=>outpp3L6(44), B=>outpp4L6(44), cin=>outpp5L6(44), S=>outpp3L4(44) ,cout=>outpp1L4(45));
FA336L6: FA port map(A=>outpp0L6(45), B=>outpp1L6(45), cin=>outpp2L6(45), S=>outpp2L4(45) ,cout=>outpp0L4(46));
FA337L6: FA port map(A=>outpp3L6(45), B=>outpp4L6(45), cin=>outpp5L6(45), S=>outpp3L4(45) ,cout=>outpp1L4(46));
FA338L6: FA port map(A=>outpp0L6(46), B=>outpp1L6(46), cin=>outpp2L6(46), S=>outpp2L4(46) ,cout=>outpp0L4(47));
FA339L6: FA port map(A=>outpp3L6(46), B=>outpp4L6(46), cin=>outpp5L6(46), S=>outpp3L4(46) ,cout=>outpp1L4(47));
FA340L6: FA port map(A=>outpp0L6(47), B=>outpp1L6(47), cin=>outpp2L6(47), S=>outpp2L4(47) ,cout=>outpp0L4(48));
FA341L6: FA port map(A=>outpp3L6(47), B=>outpp4L6(47), cin=>outpp5L6(47), S=>outpp3L4(47) ,cout=>outpp1L4(48));
FA342L6: FA port map(A=>outpp0L6(48), B=>outpp1L6(48), cin=>outpp2L6(48), S=>outpp2L4(48) ,cout=>outpp0L4(49));
FA343L6: FA port map(A=>outpp3L6(48), B=>outpp4L6(48), cin=>outpp5L6(48), S=>outpp3L4(48) ,cout=>outpp1L4(49));
FA344L6: FA port map(A=>outpp0L6(49), B=>outpp1L6(49), cin=>outpp2L6(49), S=>outpp2L4(49) ,cout=>outpp0L4(50));
FA345L6: FA port map(A=>outpp3L6(49), B=>outpp4L6(49), cin=>outpp5L6(49), S=>outpp3L4(49) ,cout=>outpp1L4(50));
FA346L6: FA port map(A=>outpp0L6(50), B=>outpp1L6(50), cin=>outpp2L6(50), S=>outpp2L4(50) ,cout=>outpp0L4(51));
FA347L6: FA port map(A=>outpp3L6(50), B=>outpp4L6(50), cin=>outpp5L6(50), S=>outpp3L4(50) ,cout=>outpp1L4(51));
FA348L6: FA port map(A=>outpp0L6(51), B=>outpp1L6(51), cin=>outpp2L6(51), S=>outpp2L4(51) ,cout=>outpp0L4(52));
FA349L6: FA port map(A=>outpp3L6(51), B=>outpp4L6(51), cin=>outpp5L6(51), S=>outpp3L4(51) ,cout=>outpp1L4(52));
FA350L6: FA port map(A=>outpp0L6(52), B=>outpp1L6(52), cin=>outpp2L6(52), S=>outpp2L4(52) ,cout=>outpp0L4(53));
FA351L6: FA port map(A=>outpp3L6(52), B=>outpp4L6(52), cin=>outpp5L6(52), S=>outpp3L4(52) ,cout=>outpp1L4(53));
FA352L6: FA port map(A=>outpp0L6(53), B=>outpp1L6(53), cin=>outpp2L6(53), S=>outpp2L4(53) ,cout=>outpp0L4(54));
FA353L6: FA port map(A=>outpp3L6(53), B=>outpp4L6(53), cin=>outpp5L6(53), S=>outpp3L4(53) ,cout=>outpp1L4(54));
FA354L6: FA port map(A=>outpp0L6(54), B=>outpp1L6(54), cin=>outpp2L6(54), S=>outpp2L4(54) ,cout=>outpp0L4(55));
FA355L6: FA port map(A=>outpp3L6(54), B=>outpp4L6(54), cin=>outpp5L6(54), S=>outpp3L4(54) ,cout=>outpp1L4(55));
FA356L6: FA port map(A=>outpp0L6(55), B=>outpp1L6(55), cin=>outpp2L6(55), S=>outpp2L4(55) ,cout=>outpp0L4(56));
FA357L6: FA port map(A=>outpp3L6(55), B=>outpp4L6(55), cin=>outpp5L6(55), S=>outpp3L4(55) ,cout=>outpp1L4(56));
FA358L6: FA port map(A=>outpp0L6(56), B=>outpp1L6(56), cin=>outpp2L6(56), S=>outpp2L4(56) ,cout=>outpp0L4(57));
FA359L6: FA port map(A=>outpp3L6(56), B=>outpp4L6(56), cin=>outpp5L6(56), S=>outpp3L4(56) ,cout=>outpp1L4(57));
FA360L6: FA port map(A=>outpp0L6(57), B=>outpp1L6(57), cin=>outpp2L6(57), S=>outpp2L4(57) ,cout=>outpp0L4(58));
FA361L6: FA port map(A=>outpp3L6(57), B=>outpp4L6(57), cin=>outpp5L6(57), S=>outpp3L4(57) ,cout=>outpp1L4(58));
HA37L6: HA port map( A=>outpp0L6(58), B=>outpp1L6(58), S=>outpp2L4(58) ,cout=>outpp0L4(59));
FA362L6: FA port map(A=>outpp2L6(58), B=>outpp3L6(58), cin=>outpp4L6(58), S=>outpp3L4(58) ,cout=>outpp1L4(59));
FA363L6: FA port map(A=>outpp0L6(59), B=>outpp1L6(59), cin=>outpp2L6(59), S=>outpp2L4(59) ,cout=>outpp0L4(60));
outpp3L4(59)<=outpp3L6(59);
HA38L6: HA port map( A=>outpp0L6(60), B=>outpp1L6(60), S=>outpp1L4(60) ,cout=>outpp0L4(61));
outpp2L4(60)<=outpp2L6(60);
outpp3L4(60)<=outpp3L6(60);
outpp1L4(61)<=outpp0L6(61);
outpp2L4(61)<=outpp1L6(61);
outpp3L4(61)<=outpp2L6(61);
outpp0L4(62)<=outpp0L6(62);
outpp1L4(62)<=outpp1L6(62);
outpp2L4(62)<=outpp2L6(62);
outpp3L4(62)<=outpp3L6(62);
outpp0L4(63)<=outpp0L6(63);
outpp1L4(63)<=outpp1L6(63);
outpp2L4(63)<=outpp2L6(63);
outpp3L4(63)<=outpp3L6(63);
outpp0L3(0)<=outpp0L4(0);
outpp1L3(0)<=outpp1L4(0);
outpp2L3(0)<=outpp2L4(0);
outpp0L3(1)<=outpp0L4(1);
outpp1L3(1)<=outpp1L4(1);
outpp2L3(1)<=outpp2L4(1);
outpp0L3(2)<=outpp0L4(2);
outpp1L3(2)<=outpp1L4(2);
outpp2L3(2)<=outpp2L4(2);
outpp0L3(3)<=outpp0L4(3);
outpp1L3(3)<=outpp1L4(3);
outpp2L3(3)<=outpp2L4(3);
HA39L4: HA port map( A=>outpp0L4(4), B=>outpp1L4(4), S=>outpp0L3(4) ,cout=>outpp0L3(5));
outpp1L3(4)<=outpp2L4(4);
outpp2L3(4)<=outpp3L4(4);
HA40L4: HA port map( A=>outpp0L4(5), B=>outpp1L4(5), S=>outpp1L3(5) ,cout=>outpp0L3(6));
outpp2L3(5)<=outpp2L4(5);
FA364L4: FA port map(A=>outpp0L4(6), B=>outpp1L4(6), cin=>outpp2L4(6), S=>outpp1L3(6) ,cout=>outpp0L3(7));
outpp2L3(6)<=outpp3L4(6);
FA365L4: FA port map(A=>outpp0L4(7), B=>outpp1L4(7), cin=>outpp2L4(7), S=>outpp1L3(7) ,cout=>outpp0L3(8));
outpp2L3(7)<=outpp3L4(7);
FA366L4: FA port map(A=>outpp0L4(8), B=>outpp1L4(8), cin=>outpp2L4(8), S=>outpp1L3(8) ,cout=>outpp0L3(9));
outpp2L3(8)<=outpp3L4(8);
FA367L4: FA port map(A=>outpp0L4(9), B=>outpp1L4(9), cin=>outpp2L4(9), S=>outpp1L3(9) ,cout=>outpp0L3(10));
outpp2L3(9)<=outpp3L4(9);
FA368L4: FA port map(A=>outpp0L4(10), B=>outpp1L4(10), cin=>outpp2L4(10), S=>outpp1L3(10) ,cout=>outpp0L3(11));
outpp2L3(10)<=outpp3L4(10);
FA369L4: FA port map(A=>outpp0L4(11), B=>outpp1L4(11), cin=>outpp2L4(11), S=>outpp1L3(11) ,cout=>outpp0L3(12));
outpp2L3(11)<=outpp3L4(11);
FA370L4: FA port map(A=>outpp0L4(12), B=>outpp1L4(12), cin=>outpp2L4(12), S=>outpp1L3(12) ,cout=>outpp0L3(13));
outpp2L3(12)<=outpp3L4(12);
FA371L4: FA port map(A=>outpp0L4(13), B=>outpp1L4(13), cin=>outpp2L4(13), S=>outpp1L3(13) ,cout=>outpp0L3(14));
outpp2L3(13)<=outpp3L4(13);
FA372L4: FA port map(A=>outpp0L4(14), B=>outpp1L4(14), cin=>outpp2L4(14), S=>outpp1L3(14) ,cout=>outpp0L3(15));
outpp2L3(14)<=outpp3L4(14);
FA373L4: FA port map(A=>outpp0L4(15), B=>outpp1L4(15), cin=>outpp2L4(15), S=>outpp1L3(15) ,cout=>outpp0L3(16));
outpp2L3(15)<=outpp3L4(15);
FA374L4: FA port map(A=>outpp0L4(16), B=>outpp1L4(16), cin=>outpp2L4(16), S=>outpp1L3(16) ,cout=>outpp0L3(17));
outpp2L3(16)<=outpp3L4(16);
FA375L4: FA port map(A=>outpp0L4(17), B=>outpp1L4(17), cin=>outpp2L4(17), S=>outpp1L3(17) ,cout=>outpp0L3(18));
outpp2L3(17)<=outpp3L4(17);
FA376L4: FA port map(A=>outpp0L4(18), B=>outpp1L4(18), cin=>outpp2L4(18), S=>outpp1L3(18) ,cout=>outpp0L3(19));
outpp2L3(18)<=outpp3L4(18);
FA377L4: FA port map(A=>outpp0L4(19), B=>outpp1L4(19), cin=>outpp2L4(19), S=>outpp1L3(19) ,cout=>outpp0L3(20));
outpp2L3(19)<=outpp3L4(19);
FA378L4: FA port map(A=>outpp0L4(20), B=>outpp1L4(20), cin=>outpp2L4(20), S=>outpp1L3(20) ,cout=>outpp0L3(21));
outpp2L3(20)<=outpp3L4(20);
FA379L4: FA port map(A=>outpp0L4(21), B=>outpp1L4(21), cin=>outpp2L4(21), S=>outpp1L3(21) ,cout=>outpp0L3(22));
outpp2L3(21)<=outpp3L4(21);
FA380L4: FA port map(A=>outpp0L4(22), B=>outpp1L4(22), cin=>outpp2L4(22), S=>outpp1L3(22) ,cout=>outpp0L3(23));
outpp2L3(22)<=outpp3L4(22);
FA381L4: FA port map(A=>outpp0L4(23), B=>outpp1L4(23), cin=>outpp2L4(23), S=>outpp1L3(23) ,cout=>outpp0L3(24));
outpp2L3(23)<=outpp3L4(23);
FA382L4: FA port map(A=>outpp0L4(24), B=>outpp1L4(24), cin=>outpp2L4(24), S=>outpp1L3(24) ,cout=>outpp0L3(25));
outpp2L3(24)<=outpp3L4(24);
FA383L4: FA port map(A=>outpp0L4(25), B=>outpp1L4(25), cin=>outpp2L4(25), S=>outpp1L3(25) ,cout=>outpp0L3(26));
outpp2L3(25)<=outpp3L4(25);
FA384L4: FA port map(A=>outpp0L4(26), B=>outpp1L4(26), cin=>outpp2L4(26), S=>outpp1L3(26) ,cout=>outpp0L3(27));
outpp2L3(26)<=outpp3L4(26);
FA385L4: FA port map(A=>outpp0L4(27), B=>outpp1L4(27), cin=>outpp2L4(27), S=>outpp1L3(27) ,cout=>outpp0L3(28));
outpp2L3(27)<=outpp3L4(27);
FA386L4: FA port map(A=>outpp0L4(28), B=>outpp1L4(28), cin=>outpp2L4(28), S=>outpp1L3(28) ,cout=>outpp0L3(29));
outpp2L3(28)<=outpp3L4(28);
FA387L4: FA port map(A=>outpp0L4(29), B=>outpp1L4(29), cin=>outpp2L4(29), S=>outpp1L3(29) ,cout=>outpp0L3(30));
outpp2L3(29)<=outpp3L4(29);
FA388L4: FA port map(A=>outpp0L4(30), B=>outpp1L4(30), cin=>outpp2L4(30), S=>outpp1L3(30) ,cout=>outpp0L3(31));
outpp2L3(30)<=outpp3L4(30);
FA389L4: FA port map(A=>outpp0L4(31), B=>outpp1L4(31), cin=>outpp2L4(31), S=>outpp1L3(31) ,cout=>outpp0L3(32));
outpp2L3(31)<=outpp3L4(31);
FA390L4: FA port map(A=>outpp0L4(32), B=>outpp1L4(32), cin=>outpp2L4(32), S=>outpp1L3(32) ,cout=>outpp0L3(33));
outpp2L3(32)<=outpp3L4(32);
FA391L4: FA port map(A=>outpp0L4(33), B=>outpp1L4(33), cin=>outpp2L4(33), S=>outpp1L3(33) ,cout=>outpp0L3(34));
outpp2L3(33)<=outpp3L4(33);
FA392L4: FA port map(A=>outpp0L4(34), B=>outpp1L4(34), cin=>outpp2L4(34), S=>outpp1L3(34) ,cout=>outpp0L3(35));
outpp2L3(34)<=outpp3L4(34);
FA393L4: FA port map(A=>outpp0L4(35), B=>outpp1L4(35), cin=>outpp2L4(35), S=>outpp1L3(35) ,cout=>outpp0L3(36));
outpp2L3(35)<=outpp3L4(35);
FA394L4: FA port map(A=>outpp0L4(36), B=>outpp1L4(36), cin=>outpp2L4(36), S=>outpp1L3(36) ,cout=>outpp0L3(37));
outpp2L3(36)<=outpp3L4(36);
FA395L4: FA port map(A=>outpp0L4(37), B=>outpp1L4(37), cin=>outpp2L4(37), S=>outpp1L3(37) ,cout=>outpp0L3(38));
outpp2L3(37)<=outpp3L4(37);
FA396L4: FA port map(A=>outpp0L4(38), B=>outpp1L4(38), cin=>outpp2L4(38), S=>outpp1L3(38) ,cout=>outpp0L3(39));
outpp2L3(38)<=outpp3L4(38);
FA397L4: FA port map(A=>outpp0L4(39), B=>outpp1L4(39), cin=>outpp2L4(39), S=>outpp1L3(39) ,cout=>outpp0L3(40));
outpp2L3(39)<=outpp3L4(39);
FA398L4: FA port map(A=>outpp0L4(40), B=>outpp1L4(40), cin=>outpp2L4(40), S=>outpp1L3(40) ,cout=>outpp0L3(41));
outpp2L3(40)<=outpp3L4(40);
FA399L4: FA port map(A=>outpp0L4(41), B=>outpp1L4(41), cin=>outpp2L4(41), S=>outpp1L3(41) ,cout=>outpp0L3(42));
outpp2L3(41)<=outpp3L4(41);
FA400L4: FA port map(A=>outpp0L4(42), B=>outpp1L4(42), cin=>outpp2L4(42), S=>outpp1L3(42) ,cout=>outpp0L3(43));
outpp2L3(42)<=outpp3L4(42);
FA401L4: FA port map(A=>outpp0L4(43), B=>outpp1L4(43), cin=>outpp2L4(43), S=>outpp1L3(43) ,cout=>outpp0L3(44));
outpp2L3(43)<=outpp3L4(43);
FA402L4: FA port map(A=>outpp0L4(44), B=>outpp1L4(44), cin=>outpp2L4(44), S=>outpp1L3(44) ,cout=>outpp0L3(45));
outpp2L3(44)<=outpp3L4(44);
FA403L4: FA port map(A=>outpp0L4(45), B=>outpp1L4(45), cin=>outpp2L4(45), S=>outpp1L3(45) ,cout=>outpp0L3(46));
outpp2L3(45)<=outpp3L4(45);
FA404L4: FA port map(A=>outpp0L4(46), B=>outpp1L4(46), cin=>outpp2L4(46), S=>outpp1L3(46) ,cout=>outpp0L3(47));
outpp2L3(46)<=outpp3L4(46);
FA405L4: FA port map(A=>outpp0L4(47), B=>outpp1L4(47), cin=>outpp2L4(47), S=>outpp1L3(47) ,cout=>outpp0L3(48));
outpp2L3(47)<=outpp3L4(47);
FA406L4: FA port map(A=>outpp0L4(48), B=>outpp1L4(48), cin=>outpp2L4(48), S=>outpp1L3(48) ,cout=>outpp0L3(49));
outpp2L3(48)<=outpp3L4(48);
FA407L4: FA port map(A=>outpp0L4(49), B=>outpp1L4(49), cin=>outpp2L4(49), S=>outpp1L3(49) ,cout=>outpp0L3(50));
outpp2L3(49)<=outpp3L4(49);
FA408L4: FA port map(A=>outpp0L4(50), B=>outpp1L4(50), cin=>outpp2L4(50), S=>outpp1L3(50) ,cout=>outpp0L3(51));
outpp2L3(50)<=outpp3L4(50);
FA409L4: FA port map(A=>outpp0L4(51), B=>outpp1L4(51), cin=>outpp2L4(51), S=>outpp1L3(51) ,cout=>outpp0L3(52));
outpp2L3(51)<=outpp3L4(51);
FA410L4: FA port map(A=>outpp0L4(52), B=>outpp1L4(52), cin=>outpp2L4(52), S=>outpp1L3(52) ,cout=>outpp0L3(53));
outpp2L3(52)<=outpp3L4(52);
FA411L4: FA port map(A=>outpp0L4(53), B=>outpp1L4(53), cin=>outpp2L4(53), S=>outpp1L3(53) ,cout=>outpp0L3(54));
outpp2L3(53)<=outpp3L4(53);
FA412L4: FA port map(A=>outpp0L4(54), B=>outpp1L4(54), cin=>outpp2L4(54), S=>outpp1L3(54) ,cout=>outpp0L3(55));
outpp2L3(54)<=outpp3L4(54);
FA413L4: FA port map(A=>outpp0L4(55), B=>outpp1L4(55), cin=>outpp2L4(55), S=>outpp1L3(55) ,cout=>outpp0L3(56));
outpp2L3(55)<=outpp3L4(55);
FA414L4: FA port map(A=>outpp0L4(56), B=>outpp1L4(56), cin=>outpp2L4(56), S=>outpp1L3(56) ,cout=>outpp0L3(57));
outpp2L3(56)<=outpp3L4(56);
FA415L4: FA port map(A=>outpp0L4(57), B=>outpp1L4(57), cin=>outpp2L4(57), S=>outpp1L3(57) ,cout=>outpp0L3(58));
outpp2L3(57)<=outpp3L4(57);
FA416L4: FA port map(A=>outpp0L4(58), B=>outpp1L4(58), cin=>outpp2L4(58), S=>outpp1L3(58) ,cout=>outpp0L3(59));
outpp2L3(58)<=outpp3L4(58);
FA417L4: FA port map(A=>outpp0L4(59), B=>outpp1L4(59), cin=>outpp2L4(59), S=>outpp1L3(59) ,cout=>outpp0L3(60));
outpp2L3(59)<=outpp3L4(59);
FA418L4: FA port map(A=>outpp0L4(60), B=>outpp1L4(60), cin=>outpp2L4(60), S=>outpp1L3(60) ,cout=>outpp0L3(61));
outpp2L3(60)<=outpp3L4(60);
FA419L4: FA port map(A=>outpp0L4(61), B=>outpp1L4(61), cin=>outpp2L4(61), S=>outpp1L3(61) ,cout=>outpp0L3(62));
outpp2L3(61)<=outpp3L4(61);
HA41L4: HA port map( A=>outpp0L4(62), B=>outpp1L4(62), S=>outpp1L3(62) ,cout=>outpp0L3(63));
outpp2L3(62)<=outpp2L4(62);
outpp1L3(63)<=outpp0L4(63);
outpp2L3(63)<=outpp1L4(63);
outpp0L2(0)<=outpp0L3(0);
outpp1L2(0)<=outpp1L3(0);
outpp0L2(1)<=outpp0L3(1);
outpp1L2(1)<=outpp1L3(1);
HA42L3: HA port map( A=>outpp0L3(2), B=>outpp1L3(2), S=>outpp0L2(2) ,cout=>outpp0L2(3));
outpp1L2(2)<=outpp2L3(2);
HA43L3: HA port map( A=>outpp0L3(3), B=>outpp1L3(3), S=>outpp1L2(3) ,cout=>outpp0L2(4));
FA420L3: FA port map(A=>outpp0L3(4), B=>outpp1L3(4), cin=>outpp2L3(4), S=>outpp1L2(4) ,cout=>outpp0L2(5));
FA421L3: FA port map(A=>outpp0L3(5), B=>outpp1L3(5), cin=>outpp2L3(5), S=>outpp1L2(5) ,cout=>outpp0L2(6));
FA422L3: FA port map(A=>outpp0L3(6), B=>outpp1L3(6), cin=>outpp2L3(6), S=>outpp1L2(6) ,cout=>outpp0L2(7));
FA423L3: FA port map(A=>outpp0L3(7), B=>outpp1L3(7), cin=>outpp2L3(7), S=>outpp1L2(7) ,cout=>outpp0L2(8));
FA424L3: FA port map(A=>outpp0L3(8), B=>outpp1L3(8), cin=>outpp2L3(8), S=>outpp1L2(8) ,cout=>outpp0L2(9));
FA425L3: FA port map(A=>outpp0L3(9), B=>outpp1L3(9), cin=>outpp2L3(9), S=>outpp1L2(9) ,cout=>outpp0L2(10));
FA426L3: FA port map(A=>outpp0L3(10), B=>outpp1L3(10), cin=>outpp2L3(10), S=>outpp1L2(10) ,cout=>outpp0L2(11));
FA427L3: FA port map(A=>outpp0L3(11), B=>outpp1L3(11), cin=>outpp2L3(11), S=>outpp1L2(11) ,cout=>outpp0L2(12));
FA428L3: FA port map(A=>outpp0L3(12), B=>outpp1L3(12), cin=>outpp2L3(12), S=>outpp1L2(12) ,cout=>outpp0L2(13));
FA429L3: FA port map(A=>outpp0L3(13), B=>outpp1L3(13), cin=>outpp2L3(13), S=>outpp1L2(13) ,cout=>outpp0L2(14));
FA430L3: FA port map(A=>outpp0L3(14), B=>outpp1L3(14), cin=>outpp2L3(14), S=>outpp1L2(14) ,cout=>outpp0L2(15));
FA431L3: FA port map(A=>outpp0L3(15), B=>outpp1L3(15), cin=>outpp2L3(15), S=>outpp1L2(15) ,cout=>outpp0L2(16));
FA432L3: FA port map(A=>outpp0L3(16), B=>outpp1L3(16), cin=>outpp2L3(16), S=>outpp1L2(16) ,cout=>outpp0L2(17));
FA433L3: FA port map(A=>outpp0L3(17), B=>outpp1L3(17), cin=>outpp2L3(17), S=>outpp1L2(17) ,cout=>outpp0L2(18));
FA434L3: FA port map(A=>outpp0L3(18), B=>outpp1L3(18), cin=>outpp2L3(18), S=>outpp1L2(18) ,cout=>outpp0L2(19));
FA435L3: FA port map(A=>outpp0L3(19), B=>outpp1L3(19), cin=>outpp2L3(19), S=>outpp1L2(19) ,cout=>outpp0L2(20));
FA436L3: FA port map(A=>outpp0L3(20), B=>outpp1L3(20), cin=>outpp2L3(20), S=>outpp1L2(20) ,cout=>outpp0L2(21));
FA437L3: FA port map(A=>outpp0L3(21), B=>outpp1L3(21), cin=>outpp2L3(21), S=>outpp1L2(21) ,cout=>outpp0L2(22));
FA438L3: FA port map(A=>outpp0L3(22), B=>outpp1L3(22), cin=>outpp2L3(22), S=>outpp1L2(22) ,cout=>outpp0L2(23));
FA439L3: FA port map(A=>outpp0L3(23), B=>outpp1L3(23), cin=>outpp2L3(23), S=>outpp1L2(23) ,cout=>outpp0L2(24));
FA440L3: FA port map(A=>outpp0L3(24), B=>outpp1L3(24), cin=>outpp2L3(24), S=>outpp1L2(24) ,cout=>outpp0L2(25));
FA441L3: FA port map(A=>outpp0L3(25), B=>outpp1L3(25), cin=>outpp2L3(25), S=>outpp1L2(25) ,cout=>outpp0L2(26));
FA442L3: FA port map(A=>outpp0L3(26), B=>outpp1L3(26), cin=>outpp2L3(26), S=>outpp1L2(26) ,cout=>outpp0L2(27));
FA443L3: FA port map(A=>outpp0L3(27), B=>outpp1L3(27), cin=>outpp2L3(27), S=>outpp1L2(27) ,cout=>outpp0L2(28));
FA444L3: FA port map(A=>outpp0L3(28), B=>outpp1L3(28), cin=>outpp2L3(28), S=>outpp1L2(28) ,cout=>outpp0L2(29));
FA445L3: FA port map(A=>outpp0L3(29), B=>outpp1L3(29), cin=>outpp2L3(29), S=>outpp1L2(29) ,cout=>outpp0L2(30));
FA446L3: FA port map(A=>outpp0L3(30), B=>outpp1L3(30), cin=>outpp2L3(30), S=>outpp1L2(30) ,cout=>outpp0L2(31));
FA447L3: FA port map(A=>outpp0L3(31), B=>outpp1L3(31), cin=>outpp2L3(31), S=>outpp1L2(31) ,cout=>outpp0L2(32));
FA448L3: FA port map(A=>outpp0L3(32), B=>outpp1L3(32), cin=>outpp2L3(32), S=>outpp1L2(32) ,cout=>outpp0L2(33));
FA449L3: FA port map(A=>outpp0L3(33), B=>outpp1L3(33), cin=>outpp2L3(33), S=>outpp1L2(33) ,cout=>outpp0L2(34));
FA450L3: FA port map(A=>outpp0L3(34), B=>outpp1L3(34), cin=>outpp2L3(34), S=>outpp1L2(34) ,cout=>outpp0L2(35));
FA451L3: FA port map(A=>outpp0L3(35), B=>outpp1L3(35), cin=>outpp2L3(35), S=>outpp1L2(35) ,cout=>outpp0L2(36));
FA452L3: FA port map(A=>outpp0L3(36), B=>outpp1L3(36), cin=>outpp2L3(36), S=>outpp1L2(36) ,cout=>outpp0L2(37));
FA453L3: FA port map(A=>outpp0L3(37), B=>outpp1L3(37), cin=>outpp2L3(37), S=>outpp1L2(37) ,cout=>outpp0L2(38));
FA454L3: FA port map(A=>outpp0L3(38), B=>outpp1L3(38), cin=>outpp2L3(38), S=>outpp1L2(38) ,cout=>outpp0L2(39));
FA455L3: FA port map(A=>outpp0L3(39), B=>outpp1L3(39), cin=>outpp2L3(39), S=>outpp1L2(39) ,cout=>outpp0L2(40));
FA456L3: FA port map(A=>outpp0L3(40), B=>outpp1L3(40), cin=>outpp2L3(40), S=>outpp1L2(40) ,cout=>outpp0L2(41));
FA457L3: FA port map(A=>outpp0L3(41), B=>outpp1L3(41), cin=>outpp2L3(41), S=>outpp1L2(41) ,cout=>outpp0L2(42));
FA458L3: FA port map(A=>outpp0L3(42), B=>outpp1L3(42), cin=>outpp2L3(42), S=>outpp1L2(42) ,cout=>outpp0L2(43));
FA459L3: FA port map(A=>outpp0L3(43), B=>outpp1L3(43), cin=>outpp2L3(43), S=>outpp1L2(43) ,cout=>outpp0L2(44));
FA460L3: FA port map(A=>outpp0L3(44), B=>outpp1L3(44), cin=>outpp2L3(44), S=>outpp1L2(44) ,cout=>outpp0L2(45));
FA461L3: FA port map(A=>outpp0L3(45), B=>outpp1L3(45), cin=>outpp2L3(45), S=>outpp1L2(45) ,cout=>outpp0L2(46));
FA462L3: FA port map(A=>outpp0L3(46), B=>outpp1L3(46), cin=>outpp2L3(46), S=>outpp1L2(46) ,cout=>outpp0L2(47));
FA463L3: FA port map(A=>outpp0L3(47), B=>outpp1L3(47), cin=>outpp2L3(47), S=>outpp1L2(47) ,cout=>outpp0L2(48));
FA464L3: FA port map(A=>outpp0L3(48), B=>outpp1L3(48), cin=>outpp2L3(48), S=>outpp1L2(48) ,cout=>outpp0L2(49));
FA465L3: FA port map(A=>outpp0L3(49), B=>outpp1L3(49), cin=>outpp2L3(49), S=>outpp1L2(49) ,cout=>outpp0L2(50));
FA466L3: FA port map(A=>outpp0L3(50), B=>outpp1L3(50), cin=>outpp2L3(50), S=>outpp1L2(50) ,cout=>outpp0L2(51));
FA467L3: FA port map(A=>outpp0L3(51), B=>outpp1L3(51), cin=>outpp2L3(51), S=>outpp1L2(51) ,cout=>outpp0L2(52));
FA468L3: FA port map(A=>outpp0L3(52), B=>outpp1L3(52), cin=>outpp2L3(52), S=>outpp1L2(52) ,cout=>outpp0L2(53));
FA469L3: FA port map(A=>outpp0L3(53), B=>outpp1L3(53), cin=>outpp2L3(53), S=>outpp1L2(53) ,cout=>outpp0L2(54));
FA470L3: FA port map(A=>outpp0L3(54), B=>outpp1L3(54), cin=>outpp2L3(54), S=>outpp1L2(54) ,cout=>outpp0L2(55));
FA471L3: FA port map(A=>outpp0L3(55), B=>outpp1L3(55), cin=>outpp2L3(55), S=>outpp1L2(55) ,cout=>outpp0L2(56));
FA472L3: FA port map(A=>outpp0L3(56), B=>outpp1L3(56), cin=>outpp2L3(56), S=>outpp1L2(56) ,cout=>outpp0L2(57));
FA473L3: FA port map(A=>outpp0L3(57), B=>outpp1L3(57), cin=>outpp2L3(57), S=>outpp1L2(57) ,cout=>outpp0L2(58));
FA474L3: FA port map(A=>outpp0L3(58), B=>outpp1L3(58), cin=>outpp2L3(58), S=>outpp1L2(58) ,cout=>outpp0L2(59));
FA475L3: FA port map(A=>outpp0L3(59), B=>outpp1L3(59), cin=>outpp2L3(59), S=>outpp1L2(59) ,cout=>outpp0L2(60));
FA476L3: FA port map(A=>outpp0L3(60), B=>outpp1L3(60), cin=>outpp2L3(60), S=>outpp1L2(60) ,cout=>outpp0L2(61));
FA477L3: FA port map(A=>outpp0L3(61), B=>outpp1L3(61), cin=>outpp2L3(61), S=>outpp1L2(61) ,cout=>outpp0L2(62));
FA478L3: FA port map(A=>outpp0L3(62), B=>outpp1L3(62), cin=>outpp2L3(62), S=>outpp1L2(62) ,cout=>outpp0L2(63));
FA479L3: FA port map(A=>outpp0L3(63), B=>outpp1L3(63), cin=>outpp2L3(63), S=>outpp1L2(63) ,cout=>outpp0L2(64));
P1<=outpp0L2(63 downto 0);
P2<=outpp1L2;
end Behavioral;
